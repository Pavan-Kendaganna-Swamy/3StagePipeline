magic
tech scmos
timestamp 1696374713
<< metal1 >>
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1013 1303 1016 1307
rect 10 1278 17 1281
rect 22 1271 25 1281
rect 82 1278 89 1281
rect 1066 1278 1073 1281
rect 1210 1278 1217 1281
rect 22 1268 33 1271
rect 70 1268 86 1271
rect 22 1262 25 1268
rect 62 1261 65 1268
rect 54 1258 65 1261
rect 118 1261 121 1271
rect 166 1268 177 1271
rect 214 1268 225 1271
rect 462 1268 470 1271
rect 542 1268 553 1271
rect 750 1268 758 1271
rect 166 1262 169 1268
rect 214 1262 217 1268
rect 114 1258 121 1261
rect 138 1258 145 1261
rect 190 1258 209 1261
rect 806 1261 809 1271
rect 822 1268 833 1271
rect 1070 1268 1078 1271
rect 1198 1268 1214 1271
rect 806 1258 825 1261
rect 922 1258 929 1261
rect 974 1258 993 1261
rect 998 1258 1014 1261
rect 1062 1258 1070 1261
rect 1218 1258 1225 1261
rect 1406 1258 1441 1261
rect 1486 1258 1502 1261
rect 974 1256 978 1258
rect 265 1248 270 1252
rect 788 1248 790 1252
rect 1406 1248 1409 1258
rect 580 1238 582 1242
rect 860 1238 862 1242
rect 1282 1238 1284 1242
rect 732 1228 734 1232
rect 421 1218 422 1222
rect 1146 1218 1148 1222
rect 488 1203 490 1207
rect 494 1203 497 1207
rect 501 1203 504 1207
rect 458 1188 459 1192
rect 756 1188 758 1192
rect 1130 1178 1131 1182
rect 906 1168 913 1171
rect 170 1158 177 1161
rect 214 1151 217 1161
rect 265 1158 270 1162
rect 1446 1158 1457 1161
rect 198 1148 217 1151
rect 438 1148 449 1151
rect 462 1148 481 1151
rect 490 1148 521 1151
rect 526 1148 542 1151
rect 594 1148 601 1151
rect 606 1148 617 1151
rect 26 1138 33 1141
rect 94 1138 113 1141
rect 206 1138 214 1141
rect 234 1138 241 1141
rect 430 1141 433 1148
rect 422 1138 433 1141
rect 446 1142 449 1148
rect 814 1148 854 1151
rect 1002 1148 1025 1151
rect 1074 1148 1081 1151
rect 1206 1151 1210 1154
rect 1182 1148 1210 1151
rect 1262 1151 1266 1154
rect 1262 1148 1273 1151
rect 774 1138 790 1141
rect 830 1138 846 1141
rect 978 1138 985 1141
rect 994 1138 1033 1141
rect 1092 1138 1121 1141
rect 1244 1138 1246 1142
rect 558 1132 561 1138
rect 394 1128 401 1131
rect 410 1128 417 1131
rect 554 1128 561 1132
rect 574 1128 593 1131
rect 830 1128 833 1138
rect 60 1118 62 1122
rect 1332 1118 1334 1122
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1013 1103 1016 1107
rect 412 1088 414 1092
rect 780 1088 782 1092
rect 818 1088 819 1092
rect 26 1078 33 1081
rect 378 1068 385 1071
rect 54 1058 65 1061
rect 430 1062 433 1071
rect 986 1068 993 1071
rect 1138 1068 1145 1071
rect 1222 1068 1241 1071
rect 1334 1071 1337 1081
rect 1318 1068 1337 1071
rect 238 1058 246 1061
rect 446 1058 454 1061
rect 950 1058 953 1068
rect 982 1058 990 1061
rect 1086 1058 1094 1061
rect 1126 1058 1150 1061
rect 1086 1056 1090 1058
rect 362 1048 369 1051
rect 1006 1048 1022 1051
rect 275 1038 278 1042
rect 532 1038 534 1042
rect 870 1038 886 1041
rect 1154 1038 1155 1042
rect 1125 1018 1126 1022
rect 488 1003 490 1007
rect 494 1003 497 1007
rect 501 1003 504 1007
rect 677 988 678 992
rect 1018 988 1019 992
rect 610 968 617 971
rect 789 968 790 972
rect 942 968 953 971
rect 1090 968 1097 971
rect 1242 968 1249 971
rect 942 962 945 968
rect 14 958 25 961
rect 750 958 758 961
rect 770 958 777 961
rect 982 958 990 961
rect 1346 958 1361 961
rect 14 948 25 951
rect 138 948 140 952
rect 22 942 25 948
rect 542 948 553 951
rect 646 948 662 951
rect 790 948 798 951
rect 802 948 817 951
rect 822 948 830 951
rect 910 951 914 954
rect 902 948 914 951
rect 1202 948 1209 951
rect 1214 948 1222 951
rect 1414 948 1425 951
rect 42 938 49 941
rect 78 938 89 941
rect 386 938 393 941
rect 634 938 641 941
rect 650 938 657 941
rect 726 938 729 948
rect 750 938 753 948
rect 902 942 905 948
rect 798 938 806 941
rect 1078 941 1081 948
rect 1078 938 1089 941
rect 1182 938 1201 941
rect 1332 938 1345 941
rect 1470 941 1473 948
rect 1470 938 1484 941
rect 46 928 49 938
rect 406 932 409 938
rect 1342 932 1345 938
rect 54 928 70 931
rect 402 928 409 932
rect 1370 918 1377 921
rect 1412 918 1414 922
rect 1466 918 1467 922
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1013 903 1016 907
rect 250 888 252 892
rect 674 888 675 892
rect 22 862 25 871
rect 46 871 49 881
rect 158 872 161 881
rect 786 878 801 881
rect 42 868 49 871
rect 70 868 81 871
rect 134 868 153 871
rect 222 868 233 871
rect 598 868 609 871
rect 702 868 713 871
rect 742 868 753 871
rect 826 868 833 871
rect 842 868 857 871
rect 874 868 881 871
rect 942 868 950 871
rect 1274 868 1281 871
rect 206 858 225 861
rect 434 858 441 861
rect 470 858 478 861
rect 710 862 713 868
rect 742 862 745 868
rect 910 858 929 861
rect 1110 858 1113 868
rect 1266 858 1289 861
rect 1398 858 1409 861
rect 470 857 474 858
rect 1398 856 1402 858
rect 14 848 25 851
rect 70 848 81 851
rect 654 848 662 851
rect 1018 848 1033 851
rect 22 842 25 848
rect 78 842 81 848
rect 1070 846 1074 848
rect 1038 838 1073 841
rect 125 818 126 822
rect 202 818 203 822
rect 1261 818 1262 822
rect 1290 818 1291 822
rect 488 803 490 807
rect 494 803 497 807
rect 501 803 504 807
rect 1306 788 1307 792
rect 602 768 609 771
rect 634 768 646 771
rect 1418 768 1433 771
rect 1062 766 1066 768
rect 1174 758 1185 761
rect 1382 758 1385 768
rect 286 756 290 758
rect 30 748 41 751
rect 38 742 41 748
rect 1382 751 1386 754
rect 1356 748 1386 751
rect 54 738 65 741
rect 110 738 118 741
rect 126 738 137 741
rect 678 741 681 748
rect 678 738 689 741
rect 790 738 798 741
rect 822 738 838 741
rect 858 738 873 741
rect 922 738 937 741
rect 950 738 974 741
rect 1042 738 1049 741
rect 1124 738 1126 742
rect 1246 738 1254 741
rect 22 728 25 738
rect 54 732 57 738
rect 382 736 386 738
rect 698 728 710 731
rect 914 728 918 732
rect 92 718 94 722
rect 1436 718 1438 722
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1013 703 1016 707
rect 212 688 214 692
rect 268 688 270 692
rect 1482 688 1484 692
rect 670 678 678 681
rect 22 671 25 678
rect 14 668 25 671
rect 178 668 185 671
rect 342 668 361 671
rect 738 668 745 671
rect 826 668 833 671
rect 974 668 982 671
rect 1070 668 1078 671
rect 1114 668 1121 671
rect 94 658 105 661
rect 158 661 161 668
rect 142 658 161 661
rect 314 658 321 661
rect 622 661 625 668
rect 614 658 625 661
rect 730 658 753 661
rect 758 658 774 661
rect 782 658 790 661
rect 846 658 854 661
rect 966 658 974 661
rect 978 658 993 661
rect 1006 658 1046 661
rect 1066 658 1089 661
rect 1106 658 1113 661
rect 598 648 606 651
rect 686 648 713 651
rect 902 651 905 658
rect 894 648 905 651
rect 1006 648 1009 658
rect 1314 648 1322 651
rect 1182 646 1186 648
rect 1318 646 1322 648
rect 802 638 809 641
rect 1182 638 1217 641
rect 1294 638 1321 641
rect 1214 628 1217 638
rect 994 618 995 622
rect 1061 618 1062 622
rect 1090 618 1091 622
rect 1492 618 1494 622
rect 488 603 490 607
rect 494 603 497 607
rect 501 603 504 607
rect 188 588 190 592
rect 706 588 707 592
rect 1238 572 1241 581
rect 1298 578 1299 582
rect 542 568 577 571
rect 1042 568 1043 572
rect 1326 568 1366 571
rect 1490 568 1491 572
rect 798 566 802 568
rect 230 558 238 561
rect 542 561 546 564
rect 542 558 550 561
rect 742 558 753 561
rect 790 558 801 561
rect 1342 558 1350 561
rect 742 552 745 558
rect 850 548 857 551
rect 1018 548 1041 551
rect 478 538 510 541
rect 566 538 569 548
rect 654 538 657 548
rect 678 538 686 541
rect 734 538 742 541
rect 814 538 822 541
rect 842 538 849 541
rect 1164 538 1177 541
rect 1398 541 1401 548
rect 1390 538 1401 541
rect 1418 538 1425 541
rect 478 536 482 538
rect 226 528 241 531
rect 262 528 281 531
rect 286 528 305 531
rect 1078 531 1081 538
rect 1174 532 1177 538
rect 1070 528 1081 531
rect 645 518 646 522
rect 757 518 758 522
rect 958 518 966 521
rect 1148 518 1150 522
rect 1322 518 1324 522
rect 1372 518 1374 522
rect 1452 518 1454 522
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1013 503 1016 507
rect 538 488 540 492
rect 346 478 353 481
rect 466 478 473 481
rect 878 478 886 481
rect 26 468 33 471
rect 14 458 30 461
rect 118 461 121 471
rect 358 471 361 478
rect 358 468 369 471
rect 438 471 441 478
rect 106 458 121 461
rect 138 458 145 461
rect 422 462 425 471
rect 438 468 446 471
rect 454 468 470 471
rect 494 468 521 471
rect 790 468 801 471
rect 854 468 865 471
rect 1046 468 1065 471
rect 1474 468 1481 471
rect 494 462 497 468
rect 390 458 398 461
rect 862 462 865 468
rect 762 458 769 461
rect 890 458 897 461
rect 982 461 985 468
rect 982 458 993 461
rect 1074 458 1089 461
rect 1406 458 1426 461
rect 1478 461 1482 464
rect 1470 458 1482 461
rect 766 448 769 458
rect 778 448 782 452
rect 958 451 961 458
rect 950 448 961 451
rect 1134 448 1142 451
rect 1398 451 1401 458
rect 1422 456 1426 458
rect 1390 448 1401 451
rect 60 438 62 442
rect 1470 438 1478 441
rect 997 418 998 422
rect 1090 418 1091 422
rect 488 403 490 407
rect 494 403 497 407
rect 501 403 504 407
rect 524 388 526 392
rect 1290 368 1329 371
rect 78 358 89 361
rect 161 358 166 362
rect 425 358 430 362
rect 986 358 990 362
rect 1002 358 1025 361
rect 1394 358 1401 361
rect 374 352 378 353
rect 30 348 38 351
rect 122 348 137 351
rect 54 338 57 348
rect 134 338 137 348
rect 750 348 766 351
rect 938 348 945 351
rect 978 348 985 351
rect 1050 348 1057 351
rect 1118 348 1126 351
rect 1182 348 1190 351
rect 1270 348 1281 351
rect 390 338 398 341
rect 490 338 497 341
rect 390 328 393 338
rect 606 332 609 342
rect 918 341 921 348
rect 1430 342 1433 351
rect 918 338 929 341
rect 1026 338 1033 341
rect 1174 338 1182 341
rect 1238 338 1246 341
rect 1346 338 1353 341
rect 1380 338 1393 341
rect 1494 338 1502 341
rect 1390 332 1393 338
rect 770 328 777 331
rect 1054 328 1065 331
rect 1150 328 1161 331
rect 1332 328 1345 331
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1013 303 1016 307
rect 694 268 702 271
rect 822 268 833 271
rect 894 271 897 281
rect 870 268 889 271
rect 894 268 913 271
rect 942 268 958 271
rect 966 268 974 271
rect 1158 268 1166 271
rect 1214 271 1217 278
rect 1214 268 1233 271
rect 1270 268 1289 271
rect 870 262 873 268
rect 1106 258 1121 261
rect 1198 258 1230 261
rect 1234 258 1241 261
rect 1246 258 1262 261
rect 1286 258 1289 268
rect 1334 258 1342 261
rect 1086 256 1090 258
rect 1086 248 1097 251
rect 203 238 206 242
rect 1366 228 1369 238
rect 488 203 490 207
rect 494 203 497 207
rect 501 203 504 207
rect 300 188 302 192
rect 1482 188 1483 192
rect 1014 168 1025 171
rect 1093 168 1094 172
rect 1266 168 1281 171
rect 1324 168 1326 172
rect 726 166 730 168
rect 1022 162 1025 168
rect 38 148 54 151
rect 358 148 366 151
rect 482 148 489 151
rect 718 148 737 151
rect 798 151 801 158
rect 798 148 809 151
rect 990 148 1017 151
rect 1438 151 1442 153
rect 734 142 737 148
rect 446 138 454 141
rect 462 138 481 141
rect 742 138 761 141
rect 822 141 825 148
rect 814 138 825 141
rect 886 138 897 141
rect 974 141 977 148
rect 1438 148 1449 151
rect 1474 148 1481 151
rect 964 138 977 141
rect 1154 138 1161 141
rect 1284 138 1297 141
rect 478 128 481 138
rect 758 128 761 138
rect 906 128 913 131
rect 1146 128 1153 131
rect 1180 128 1206 131
rect 138 118 140 122
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1013 103 1016 107
rect 36 88 38 92
rect 148 88 150 92
rect 252 88 254 92
rect 370 88 372 92
rect 494 88 510 91
rect 214 71 217 81
rect 170 68 177 71
rect 198 68 209 71
rect 214 68 222 71
rect 846 68 858 71
rect 910 68 913 78
rect 254 58 281 61
rect 294 58 310 61
rect 326 61 329 68
rect 326 58 337 61
rect 630 58 642 61
rect 750 58 762 61
rect 66 48 73 51
rect 278 48 281 58
rect 638 57 642 58
rect 758 57 762 58
rect 942 58 953 61
rect 1078 58 1089 61
rect 1198 58 1209 61
rect 1318 58 1329 61
rect 1438 58 1449 61
rect 942 57 946 58
rect 1078 57 1082 58
rect 1198 57 1202 58
rect 1318 57 1322 58
rect 1438 57 1442 58
rect 488 3 490 7
rect 494 3 497 7
rect 501 3 504 7
<< m2contact >>
rect 1002 1303 1006 1307
rect 1009 1303 1013 1307
rect 294 1288 298 1292
rect 1070 1288 1074 1292
rect 6 1278 10 1282
rect 62 1278 66 1282
rect 78 1278 82 1282
rect 214 1278 218 1282
rect 230 1278 234 1282
rect 430 1278 434 1282
rect 486 1278 490 1282
rect 534 1278 538 1282
rect 1062 1278 1066 1282
rect 1206 1278 1210 1282
rect 1350 1278 1354 1282
rect 1470 1278 1474 1282
rect 62 1268 66 1272
rect 86 1268 90 1272
rect 102 1268 106 1272
rect 6 1258 10 1262
rect 22 1258 26 1262
rect 38 1258 42 1262
rect 78 1258 82 1262
rect 94 1258 98 1262
rect 110 1258 114 1262
rect 198 1268 202 1272
rect 238 1268 242 1272
rect 286 1268 290 1272
rect 310 1268 314 1272
rect 350 1268 354 1272
rect 470 1268 474 1272
rect 510 1268 514 1272
rect 598 1268 602 1272
rect 614 1268 618 1272
rect 702 1268 706 1272
rect 758 1268 762 1272
rect 134 1258 138 1262
rect 166 1258 170 1262
rect 214 1258 218 1262
rect 342 1259 346 1263
rect 374 1258 378 1262
rect 414 1258 418 1262
rect 454 1258 458 1262
rect 470 1258 474 1262
rect 630 1259 634 1263
rect 662 1258 666 1262
rect 814 1268 818 1272
rect 878 1268 882 1272
rect 942 1268 946 1272
rect 1006 1268 1010 1272
rect 1078 1268 1082 1272
rect 1094 1268 1098 1272
rect 1126 1268 1130 1272
rect 1174 1268 1178 1272
rect 1190 1268 1194 1272
rect 1214 1268 1218 1272
rect 1262 1268 1266 1272
rect 1310 1268 1314 1272
rect 1358 1268 1362 1272
rect 1366 1268 1370 1272
rect 1382 1268 1386 1272
rect 1414 1268 1418 1272
rect 1462 1268 1466 1272
rect 894 1258 898 1262
rect 918 1258 922 1262
rect 934 1258 938 1262
rect 966 1258 970 1262
rect 1014 1258 1018 1262
rect 1070 1258 1074 1262
rect 1102 1258 1106 1262
rect 1110 1258 1114 1262
rect 1182 1258 1186 1262
rect 1214 1258 1218 1262
rect 1238 1258 1242 1262
rect 1326 1258 1330 1262
rect 1374 1258 1378 1262
rect 1390 1258 1394 1262
rect 1398 1258 1402 1262
rect 1502 1258 1506 1262
rect 174 1248 178 1252
rect 270 1248 274 1252
rect 294 1248 298 1252
rect 438 1248 442 1252
rect 478 1248 482 1252
rect 526 1248 530 1252
rect 790 1248 794 1252
rect 886 1248 890 1252
rect 918 1248 922 1252
rect 982 1248 986 1252
rect 1118 1248 1122 1252
rect 1230 1248 1234 1252
rect 1318 1248 1322 1252
rect 582 1238 586 1242
rect 862 1238 866 1242
rect 902 1238 906 1242
rect 958 1238 962 1242
rect 1246 1238 1250 1242
rect 1278 1238 1282 1242
rect 1334 1238 1338 1242
rect 734 1228 738 1232
rect 1342 1228 1346 1232
rect 406 1218 410 1222
rect 422 1218 426 1222
rect 518 1218 522 1222
rect 694 1218 698 1222
rect 910 1218 914 1222
rect 966 1218 970 1222
rect 1142 1218 1146 1222
rect 1254 1218 1258 1222
rect 1486 1218 1490 1222
rect 490 1203 494 1207
rect 497 1203 501 1207
rect 454 1188 458 1192
rect 758 1188 762 1192
rect 790 1188 794 1192
rect 902 1188 906 1192
rect 958 1188 962 1192
rect 1046 1188 1050 1192
rect 1230 1188 1234 1192
rect 934 1178 938 1182
rect 1126 1178 1130 1182
rect 1438 1178 1442 1182
rect 902 1168 906 1172
rect 950 1168 954 1172
rect 1222 1168 1226 1172
rect 1246 1168 1250 1172
rect 1358 1168 1362 1172
rect 1366 1168 1370 1172
rect 1430 1168 1434 1172
rect 22 1158 26 1162
rect 166 1158 170 1162
rect 206 1158 210 1162
rect 102 1148 106 1152
rect 190 1148 194 1152
rect 270 1158 274 1162
rect 534 1158 538 1162
rect 558 1158 562 1162
rect 870 1158 874 1162
rect 894 1158 898 1162
rect 966 1158 970 1162
rect 1142 1158 1146 1162
rect 1206 1158 1210 1162
rect 1262 1158 1266 1162
rect 1382 1158 1386 1162
rect 318 1147 322 1151
rect 350 1148 354 1152
rect 390 1148 394 1152
rect 430 1148 434 1152
rect 486 1148 490 1152
rect 542 1148 546 1152
rect 582 1148 586 1152
rect 590 1148 594 1152
rect 6 1138 10 1142
rect 22 1138 26 1142
rect 78 1138 82 1142
rect 158 1138 162 1142
rect 182 1138 186 1142
rect 214 1138 218 1142
rect 230 1138 234 1142
rect 286 1138 290 1142
rect 654 1147 658 1151
rect 854 1148 858 1152
rect 862 1148 866 1152
rect 902 1148 906 1152
rect 958 1148 962 1152
rect 998 1148 1002 1152
rect 1070 1148 1074 1152
rect 1126 1148 1130 1152
rect 1214 1148 1218 1152
rect 1254 1148 1258 1152
rect 1374 1148 1378 1152
rect 1390 1148 1394 1152
rect 1438 1148 1442 1152
rect 1494 1148 1498 1152
rect 446 1138 450 1142
rect 510 1138 514 1142
rect 542 1138 546 1142
rect 558 1138 562 1142
rect 662 1138 666 1142
rect 790 1138 794 1142
rect 814 1138 818 1142
rect 846 1138 850 1142
rect 974 1138 978 1142
rect 990 1138 994 1142
rect 1070 1138 1074 1142
rect 1078 1138 1082 1142
rect 1150 1138 1154 1142
rect 1198 1138 1202 1142
rect 1246 1138 1250 1142
rect 1278 1138 1282 1142
rect 1302 1138 1306 1142
rect 1350 1138 1354 1142
rect 1398 1138 1402 1142
rect 1486 1138 1490 1142
rect 86 1128 90 1132
rect 166 1128 170 1132
rect 390 1128 394 1132
rect 406 1128 410 1132
rect 430 1128 434 1132
rect 446 1128 450 1132
rect 470 1128 474 1132
rect 566 1128 570 1132
rect 622 1128 626 1132
rect 886 1128 890 1132
rect 926 1128 930 1132
rect 974 1128 978 1132
rect 1046 1128 1050 1132
rect 1062 1128 1066 1132
rect 1294 1128 1298 1132
rect 1414 1128 1418 1132
rect 1462 1128 1466 1132
rect 1470 1128 1474 1132
rect 22 1118 26 1122
rect 62 1118 66 1122
rect 134 1118 138 1122
rect 214 1118 218 1122
rect 382 1118 386 1122
rect 718 1118 722 1122
rect 878 1118 882 1122
rect 1286 1118 1290 1122
rect 1334 1118 1338 1122
rect 1406 1118 1410 1122
rect 1478 1118 1482 1122
rect 1002 1103 1006 1107
rect 1009 1103 1013 1107
rect 14 1088 18 1092
rect 70 1088 74 1092
rect 198 1088 202 1092
rect 294 1088 298 1092
rect 414 1088 418 1092
rect 782 1088 786 1092
rect 814 1088 818 1092
rect 846 1088 850 1092
rect 902 1088 906 1092
rect 934 1088 938 1092
rect 1342 1088 1346 1092
rect 1502 1088 1506 1092
rect 6 1078 10 1082
rect 22 1078 26 1082
rect 38 1078 42 1082
rect 46 1078 50 1082
rect 78 1078 82 1082
rect 438 1078 442 1082
rect 854 1078 858 1082
rect 926 1078 930 1082
rect 982 1078 986 1082
rect 1094 1078 1098 1082
rect 1230 1078 1234 1082
rect 1326 1078 1330 1082
rect 86 1068 90 1072
rect 230 1068 234 1072
rect 302 1068 306 1072
rect 350 1068 354 1072
rect 358 1068 362 1072
rect 374 1068 378 1072
rect 22 1058 26 1062
rect 134 1059 138 1063
rect 462 1068 466 1072
rect 478 1068 482 1072
rect 502 1068 506 1072
rect 550 1068 554 1072
rect 662 1068 666 1072
rect 750 1068 754 1072
rect 798 1068 802 1072
rect 806 1068 810 1072
rect 838 1068 842 1072
rect 942 1068 946 1072
rect 950 1068 954 1072
rect 966 1068 970 1072
rect 982 1068 986 1072
rect 1070 1068 1074 1072
rect 1134 1068 1138 1072
rect 1214 1068 1218 1072
rect 1254 1068 1258 1072
rect 1310 1068 1314 1072
rect 1510 1078 1514 1082
rect 1350 1068 1354 1072
rect 1366 1068 1370 1072
rect 1414 1068 1418 1072
rect 1422 1068 1426 1072
rect 1494 1068 1498 1072
rect 166 1058 170 1062
rect 246 1058 250 1062
rect 430 1058 434 1062
rect 454 1058 458 1062
rect 470 1058 474 1062
rect 582 1059 586 1063
rect 614 1058 618 1062
rect 686 1058 690 1062
rect 830 1058 834 1062
rect 878 1058 882 1062
rect 910 1058 914 1062
rect 958 1058 962 1062
rect 990 1058 994 1062
rect 1046 1058 1050 1062
rect 1078 1058 1082 1062
rect 1094 1058 1098 1062
rect 1150 1058 1154 1062
rect 1190 1058 1194 1062
rect 1206 1058 1210 1062
rect 1246 1058 1250 1062
rect 1286 1058 1290 1062
rect 1302 1058 1306 1062
rect 1358 1058 1362 1062
rect 1382 1058 1386 1062
rect 1430 1058 1434 1062
rect 1438 1058 1442 1062
rect 1470 1058 1474 1062
rect 1486 1058 1490 1062
rect 102 1048 106 1052
rect 358 1048 362 1052
rect 374 1048 378 1052
rect 454 1048 458 1052
rect 822 1048 826 1052
rect 886 1048 890 1052
rect 918 1048 922 1052
rect 1022 1048 1026 1052
rect 1054 1048 1058 1052
rect 1086 1048 1090 1052
rect 1110 1048 1114 1052
rect 1166 1048 1170 1052
rect 1198 1048 1202 1052
rect 1262 1048 1266 1052
rect 1294 1048 1298 1052
rect 1446 1048 1450 1052
rect 1478 1048 1482 1052
rect 278 1038 282 1042
rect 534 1038 538 1042
rect 886 1038 890 1042
rect 902 1038 906 1042
rect 1038 1038 1042 1042
rect 1070 1038 1074 1042
rect 1150 1038 1154 1042
rect 1182 1038 1186 1042
rect 1278 1038 1282 1042
rect 1462 1038 1466 1042
rect 878 1028 882 1032
rect 1046 1028 1050 1032
rect 1102 1028 1106 1032
rect 1190 1028 1194 1032
rect 94 1018 98 1022
rect 326 1018 330 1022
rect 646 1018 650 1022
rect 742 1018 746 1022
rect 998 1018 1002 1022
rect 1126 1018 1130 1022
rect 1286 1018 1290 1022
rect 1470 1018 1474 1022
rect 490 1003 494 1007
rect 497 1003 501 1007
rect 358 988 362 992
rect 542 988 546 992
rect 678 988 682 992
rect 846 988 850 992
rect 870 988 874 992
rect 894 988 898 992
rect 918 988 922 992
rect 974 988 978 992
rect 1014 988 1018 992
rect 1118 988 1122 992
rect 1278 988 1282 992
rect 262 968 266 972
rect 606 968 610 972
rect 790 968 794 972
rect 926 968 930 972
rect 1086 968 1090 972
rect 1126 968 1130 972
rect 1238 968 1242 972
rect 1270 968 1274 972
rect 1302 968 1306 972
rect 1334 968 1338 972
rect 1374 968 1378 972
rect 1406 968 1410 972
rect 1486 968 1490 972
rect 406 958 410 962
rect 598 958 602 962
rect 718 958 722 962
rect 758 958 762 962
rect 766 958 770 962
rect 830 958 834 962
rect 854 958 858 962
rect 878 958 882 962
rect 886 958 890 962
rect 942 958 946 962
rect 958 958 962 962
rect 990 958 994 962
rect 1102 958 1106 962
rect 1110 958 1114 962
rect 1222 958 1226 962
rect 1230 958 1234 962
rect 1254 958 1258 962
rect 1286 958 1290 962
rect 1318 958 1322 962
rect 1342 958 1346 962
rect 1390 958 1394 962
rect 1470 958 1474 962
rect 1502 958 1506 962
rect 62 948 66 952
rect 134 948 138 952
rect 198 947 202 951
rect 230 948 234 952
rect 302 948 306 952
rect 382 948 386 952
rect 438 947 442 951
rect 470 948 474 952
rect 590 948 594 952
rect 606 948 610 952
rect 662 948 666 952
rect 678 948 682 952
rect 702 948 706 952
rect 726 948 730 952
rect 734 948 738 952
rect 750 948 754 952
rect 798 948 802 952
rect 830 948 834 952
rect 918 948 922 952
rect 1014 948 1018 952
rect 1030 948 1034 952
rect 1046 948 1050 952
rect 1078 948 1082 952
rect 1118 948 1122 952
rect 1142 948 1146 952
rect 1158 948 1162 952
rect 1174 948 1178 952
rect 1198 948 1202 952
rect 1222 948 1226 952
rect 1238 948 1242 952
rect 1278 948 1282 952
rect 1310 948 1314 952
rect 1342 948 1346 952
rect 1366 948 1370 952
rect 1398 948 1402 952
rect 1470 948 1474 952
rect 1494 948 1498 952
rect 22 938 26 942
rect 30 938 34 942
rect 38 938 42 942
rect 94 940 98 944
rect 118 938 122 942
rect 166 938 170 942
rect 206 938 210 942
rect 278 938 282 942
rect 310 938 314 942
rect 382 938 386 942
rect 406 938 410 942
rect 582 938 586 942
rect 630 938 634 942
rect 646 938 650 942
rect 686 938 690 942
rect 694 938 698 942
rect 806 938 810 942
rect 838 938 842 942
rect 862 938 866 942
rect 902 938 906 942
rect 942 938 946 942
rect 966 938 970 942
rect 1006 938 1010 942
rect 1038 938 1042 942
rect 1054 938 1058 942
rect 1070 938 1074 942
rect 1150 938 1154 942
rect 1430 938 1434 942
rect 1454 938 1458 942
rect 6 928 10 932
rect 70 928 74 932
rect 366 928 370 932
rect 526 928 530 932
rect 558 928 562 932
rect 566 928 570 932
rect 630 928 634 932
rect 766 928 770 932
rect 1062 928 1066 932
rect 1166 928 1170 932
rect 1190 928 1194 932
rect 1342 928 1346 932
rect 1446 928 1450 932
rect 78 918 82 922
rect 110 918 114 922
rect 374 918 378 922
rect 502 918 506 922
rect 574 918 578 922
rect 614 918 618 922
rect 718 918 722 922
rect 1302 918 1306 922
rect 1366 918 1370 922
rect 1414 918 1418 922
rect 1438 918 1442 922
rect 1462 918 1466 922
rect 1002 903 1006 907
rect 1009 903 1013 907
rect 102 888 106 892
rect 166 888 170 892
rect 246 888 250 892
rect 374 888 378 892
rect 630 888 634 892
rect 654 888 658 892
rect 670 888 674 892
rect 686 888 690 892
rect 726 888 730 892
rect 766 888 770 892
rect 806 888 810 892
rect 862 888 866 892
rect 1030 888 1034 892
rect 1206 888 1210 892
rect 1318 888 1322 892
rect 1422 888 1426 892
rect 6 878 10 882
rect 38 868 42 872
rect 142 878 146 882
rect 150 878 154 882
rect 190 878 194 882
rect 310 878 314 882
rect 590 878 594 882
rect 838 878 842 882
rect 870 878 874 882
rect 902 878 906 882
rect 1110 878 1114 882
rect 1174 878 1178 882
rect 1222 878 1226 882
rect 1310 878 1314 882
rect 1430 878 1434 882
rect 54 868 58 872
rect 158 868 162 872
rect 174 868 178 872
rect 214 868 218 872
rect 278 868 282 872
rect 502 868 506 872
rect 638 868 642 872
rect 662 868 666 872
rect 718 868 722 872
rect 734 868 738 872
rect 774 868 778 872
rect 814 868 818 872
rect 822 868 826 872
rect 838 868 842 872
rect 870 868 874 872
rect 918 868 922 872
rect 950 868 954 872
rect 958 868 962 872
rect 974 868 978 872
rect 990 868 994 872
rect 1046 868 1050 872
rect 1094 868 1098 872
rect 1110 868 1114 872
rect 1158 868 1162 872
rect 1166 868 1170 872
rect 1182 868 1186 872
rect 1214 868 1218 872
rect 1270 868 1274 872
rect 1326 868 1330 872
rect 1414 868 1418 872
rect 22 858 26 862
rect 86 858 90 862
rect 126 858 130 862
rect 182 858 186 862
rect 310 859 314 863
rect 406 859 410 863
rect 430 858 434 862
rect 478 858 482 862
rect 518 859 522 863
rect 614 858 618 862
rect 710 858 714 862
rect 742 858 746 862
rect 822 858 826 862
rect 846 858 850 862
rect 950 858 954 862
rect 982 858 986 862
rect 1062 858 1066 862
rect 1086 858 1090 862
rect 1126 858 1130 862
rect 1150 858 1154 862
rect 1190 858 1194 862
rect 1206 858 1210 862
rect 1238 858 1242 862
rect 1262 858 1266 862
rect 1334 858 1338 862
rect 1358 858 1362 862
rect 1390 858 1394 862
rect 1446 858 1450 862
rect 1478 858 1482 862
rect 38 848 42 852
rect 110 848 114 852
rect 662 848 666 852
rect 678 848 682 852
rect 686 848 690 852
rect 766 848 770 852
rect 790 848 794 852
rect 894 848 898 852
rect 942 848 946 852
rect 1006 848 1010 852
rect 1014 848 1018 852
rect 1054 848 1058 852
rect 1070 848 1074 852
rect 1118 848 1122 852
rect 1246 848 1250 852
rect 1302 848 1306 852
rect 1366 848 1370 852
rect 1398 848 1402 852
rect 1438 848 1442 852
rect 1470 848 1474 852
rect 22 838 26 842
rect 30 838 34 842
rect 78 838 82 842
rect 1134 838 1138 842
rect 1238 838 1242 842
rect 1350 838 1354 842
rect 1382 838 1386 842
rect 1454 838 1458 842
rect 1486 838 1490 842
rect 886 828 890 832
rect 126 818 130 822
rect 198 818 202 822
rect 582 818 586 822
rect 958 818 962 822
rect 998 818 1002 822
rect 1078 818 1082 822
rect 1126 818 1130 822
rect 1262 818 1266 822
rect 1286 818 1290 822
rect 1358 818 1362 822
rect 1390 818 1394 822
rect 1430 818 1434 822
rect 1446 818 1450 822
rect 1478 818 1482 822
rect 490 803 494 807
rect 497 803 501 807
rect 758 788 762 792
rect 1182 788 1186 792
rect 1302 788 1306 792
rect 1502 788 1506 792
rect 638 778 642 782
rect 1390 778 1394 782
rect 590 768 594 772
rect 598 768 602 772
rect 630 768 634 772
rect 646 768 650 772
rect 1062 768 1066 772
rect 1126 768 1130 772
rect 1158 768 1162 772
rect 1214 768 1218 772
rect 1278 768 1282 772
rect 1382 768 1386 772
rect 1398 768 1402 772
rect 1414 768 1418 772
rect 1454 768 1458 772
rect 158 758 162 762
rect 286 758 290 762
rect 614 758 618 762
rect 646 758 650 762
rect 702 758 706 762
rect 854 758 858 762
rect 918 758 922 762
rect 1110 758 1114 762
rect 1142 758 1146 762
rect 1198 758 1202 762
rect 1262 758 1266 762
rect 1286 758 1290 762
rect 1318 758 1322 762
rect 1414 758 1418 762
rect 1470 758 1474 762
rect 54 748 58 752
rect 142 748 146 752
rect 150 748 154 752
rect 190 748 194 752
rect 222 747 226 751
rect 318 747 322 751
rect 350 748 354 752
rect 414 747 418 751
rect 526 747 530 751
rect 638 748 642 752
rect 678 748 682 752
rect 718 748 722 752
rect 734 748 738 752
rect 742 748 746 752
rect 774 748 778 752
rect 806 748 810 752
rect 862 748 866 752
rect 894 748 898 752
rect 926 748 930 752
rect 958 748 962 752
rect 966 748 970 752
rect 1014 748 1018 752
rect 1086 748 1090 752
rect 1134 748 1138 752
rect 1166 748 1170 752
rect 1206 748 1210 752
rect 1230 748 1234 752
rect 1270 748 1274 752
rect 1302 748 1306 752
rect 1390 748 1394 752
rect 1422 748 1426 752
rect 1462 748 1466 752
rect 1478 748 1482 752
rect 22 738 26 742
rect 38 738 42 742
rect 118 738 122 742
rect 182 738 186 742
rect 206 738 210 742
rect 382 738 386 742
rect 430 738 434 742
rect 598 738 602 742
rect 670 738 674 742
rect 726 738 730 742
rect 798 738 802 742
rect 838 738 842 742
rect 854 738 858 742
rect 886 738 890 742
rect 902 738 906 742
rect 918 738 922 742
rect 974 738 978 742
rect 1022 738 1026 742
rect 1038 738 1042 742
rect 1094 738 1098 742
rect 1126 738 1130 742
rect 1190 738 1194 742
rect 1238 738 1242 742
rect 1254 738 1258 742
rect 1294 738 1298 742
rect 1326 738 1330 742
rect 1374 738 1378 742
rect 1486 738 1490 742
rect 6 728 10 732
rect 38 728 42 732
rect 54 728 58 732
rect 118 728 122 732
rect 166 728 170 732
rect 526 728 530 732
rect 654 728 658 732
rect 710 728 714 732
rect 918 728 922 732
rect 990 728 994 732
rect 1038 728 1042 732
rect 1054 728 1058 732
rect 1070 728 1074 732
rect 1254 728 1258 732
rect 1502 728 1506 732
rect 14 718 18 722
rect 46 718 50 722
rect 94 718 98 722
rect 174 718 178 722
rect 478 718 482 722
rect 662 718 666 722
rect 758 718 762 722
rect 854 718 858 722
rect 878 718 882 722
rect 942 718 946 722
rect 982 718 986 722
rect 1030 718 1034 722
rect 1078 718 1082 722
rect 1110 718 1114 722
rect 1158 718 1162 722
rect 1214 718 1218 722
rect 1438 718 1442 722
rect 1454 718 1458 722
rect 1002 703 1006 707
rect 1009 703 1013 707
rect 158 688 162 692
rect 214 688 218 692
rect 270 688 274 692
rect 574 688 578 692
rect 598 688 602 692
rect 870 688 874 692
rect 1126 688 1130 692
rect 1382 688 1386 692
rect 1478 688 1482 692
rect 6 678 10 682
rect 22 678 26 682
rect 86 678 90 682
rect 126 678 130 682
rect 150 678 154 682
rect 350 678 354 682
rect 678 678 682 682
rect 694 678 698 682
rect 934 678 938 682
rect 1134 678 1138 682
rect 1254 678 1258 682
rect 1262 678 1266 682
rect 1390 678 1394 682
rect 30 668 34 672
rect 110 668 114 672
rect 158 668 162 672
rect 174 668 178 672
rect 230 668 234 672
rect 238 668 242 672
rect 286 668 290 672
rect 294 668 298 672
rect 494 668 498 672
rect 526 668 530 672
rect 582 668 586 672
rect 606 668 610 672
rect 622 668 626 672
rect 734 668 738 672
rect 774 668 778 672
rect 798 668 802 672
rect 822 668 826 672
rect 902 668 906 672
rect 910 668 914 672
rect 942 668 946 672
rect 982 668 986 672
rect 1030 668 1034 672
rect 1078 668 1082 672
rect 1110 668 1114 672
rect 1246 668 1250 672
rect 1374 668 1378 672
rect 1462 668 1466 672
rect 1510 668 1514 672
rect 22 658 26 662
rect 134 658 138 662
rect 310 658 314 662
rect 366 658 370 662
rect 398 659 402 663
rect 430 658 434 662
rect 510 659 514 663
rect 646 658 650 662
rect 678 658 682 662
rect 718 658 722 662
rect 726 658 730 662
rect 774 658 778 662
rect 790 658 794 662
rect 854 658 858 662
rect 902 658 906 662
rect 918 658 922 662
rect 934 658 938 662
rect 958 658 962 662
rect 974 658 978 662
rect 1046 658 1050 662
rect 1062 658 1066 662
rect 1102 658 1106 662
rect 1150 658 1154 662
rect 1190 658 1194 662
rect 1214 658 1218 662
rect 1238 658 1242 662
rect 1278 658 1282 662
rect 1310 658 1314 662
rect 1342 658 1346 662
rect 1366 658 1370 662
rect 1414 658 1418 662
rect 1446 658 1450 662
rect 158 648 162 652
rect 606 648 610 652
rect 622 648 626 652
rect 654 648 658 652
rect 766 648 770 652
rect 790 648 794 652
rect 814 648 818 652
rect 886 648 890 652
rect 950 648 954 652
rect 1046 648 1050 652
rect 1102 648 1106 652
rect 1142 648 1146 652
rect 1182 648 1186 652
rect 1198 648 1202 652
rect 1206 648 1210 652
rect 1270 648 1274 652
rect 1302 648 1306 652
rect 1310 648 1314 652
rect 1334 648 1338 652
rect 1422 648 1426 652
rect 1454 648 1458 652
rect 638 638 642 642
rect 670 638 674 642
rect 798 638 802 642
rect 1158 638 1162 642
rect 1222 638 1226 642
rect 1286 638 1290 642
rect 1350 638 1354 642
rect 1406 638 1410 642
rect 1438 638 1442 642
rect 646 628 650 632
rect 54 618 58 622
rect 126 618 130 622
rect 462 618 466 622
rect 990 618 994 622
rect 1062 618 1066 622
rect 1086 618 1090 622
rect 1150 618 1154 622
rect 1174 618 1178 622
rect 1310 618 1314 622
rect 1342 618 1346 622
rect 1398 618 1402 622
rect 1430 618 1434 622
rect 1494 618 1498 622
rect 490 603 494 607
rect 497 603 501 607
rect 190 588 194 592
rect 310 588 314 592
rect 478 588 482 592
rect 526 588 530 592
rect 550 588 554 592
rect 702 588 706 592
rect 1294 578 1298 582
rect 798 568 802 572
rect 934 568 938 572
rect 958 568 962 572
rect 1038 568 1042 572
rect 1070 568 1074 572
rect 1142 568 1146 572
rect 1166 568 1170 572
rect 1230 568 1234 572
rect 1238 568 1242 572
rect 1366 568 1370 572
rect 1486 568 1490 572
rect 238 558 242 562
rect 246 558 250 562
rect 550 558 554 562
rect 558 558 562 562
rect 582 558 586 562
rect 606 558 610 562
rect 630 558 634 562
rect 638 558 642 562
rect 718 558 722 562
rect 918 558 922 562
rect 942 558 946 562
rect 974 558 978 562
rect 1054 558 1058 562
rect 1086 558 1090 562
rect 1126 558 1130 562
rect 1182 558 1186 562
rect 1246 558 1250 562
rect 1310 558 1314 562
rect 1350 558 1354 562
rect 1398 558 1402 562
rect 1502 558 1506 562
rect 38 548 42 552
rect 86 547 90 551
rect 118 548 122 552
rect 270 548 274 552
rect 294 548 298 552
rect 326 548 330 552
rect 422 548 426 552
rect 502 548 506 552
rect 550 548 554 552
rect 566 548 570 552
rect 654 548 658 552
rect 662 548 666 552
rect 702 548 706 552
rect 742 548 746 552
rect 838 548 842 552
rect 846 548 850 552
rect 870 548 874 552
rect 910 548 914 552
rect 926 548 930 552
rect 966 548 970 552
rect 982 548 986 552
rect 1014 548 1018 552
rect 1078 548 1082 552
rect 1094 548 1098 552
rect 1134 548 1138 552
rect 1174 548 1178 552
rect 1190 548 1194 552
rect 1238 548 1242 552
rect 1278 548 1282 552
rect 1294 548 1298 552
rect 1334 548 1338 552
rect 1358 548 1362 552
rect 1398 548 1402 552
rect 1486 548 1490 552
rect 54 538 58 542
rect 206 538 210 542
rect 214 538 218 542
rect 382 538 386 542
rect 398 538 402 542
rect 430 538 434 542
rect 510 538 514 542
rect 590 538 594 542
rect 614 538 618 542
rect 686 538 690 542
rect 694 538 698 542
rect 726 538 730 542
rect 742 538 746 542
rect 766 538 770 542
rect 774 538 778 542
rect 822 538 826 542
rect 838 538 842 542
rect 878 538 882 542
rect 902 538 906 542
rect 990 538 994 542
rect 1030 538 1034 542
rect 1078 538 1082 542
rect 1102 538 1106 542
rect 1198 538 1202 542
rect 1270 538 1274 542
rect 1286 538 1290 542
rect 1382 538 1386 542
rect 1414 538 1418 542
rect 1470 538 1474 542
rect 1478 538 1482 542
rect 254 528 258 532
rect 526 528 530 532
rect 806 528 810 532
rect 822 528 826 532
rect 870 528 874 532
rect 886 528 890 532
rect 1006 528 1010 532
rect 1118 528 1122 532
rect 1174 528 1178 532
rect 1214 528 1218 532
rect 1254 528 1258 532
rect 1262 528 1266 532
rect 150 518 154 522
rect 582 518 586 522
rect 606 518 610 522
rect 630 518 634 522
rect 646 518 650 522
rect 758 518 762 522
rect 790 518 794 522
rect 830 518 834 522
rect 894 518 898 522
rect 966 518 970 522
rect 998 518 1002 522
rect 1110 518 1114 522
rect 1150 518 1154 522
rect 1206 518 1210 522
rect 1318 518 1322 522
rect 1374 518 1378 522
rect 1406 518 1410 522
rect 1454 518 1458 522
rect 1002 503 1006 507
rect 1009 503 1013 507
rect 86 488 90 492
rect 262 488 266 492
rect 478 488 482 492
rect 534 488 538 492
rect 662 488 666 492
rect 814 488 818 492
rect 870 488 874 492
rect 926 488 930 492
rect 1038 488 1042 492
rect 1166 488 1170 492
rect 1230 488 1234 492
rect 1342 488 1346 492
rect 342 478 346 482
rect 358 478 362 482
rect 430 478 434 482
rect 438 478 442 482
rect 446 478 450 482
rect 462 478 466 482
rect 742 478 746 482
rect 806 478 810 482
rect 862 478 866 482
rect 886 478 890 482
rect 1006 478 1010 482
rect 1030 478 1034 482
rect 1070 478 1074 482
rect 1142 478 1146 482
rect 1158 478 1162 482
rect 1262 478 1266 482
rect 1334 478 1338 482
rect 1366 478 1370 482
rect 1454 478 1458 482
rect 6 468 10 472
rect 22 468 26 472
rect 110 468 114 472
rect 30 458 34 462
rect 102 458 106 462
rect 166 468 170 472
rect 182 468 186 472
rect 334 468 338 472
rect 398 468 402 472
rect 134 458 138 462
rect 198 459 202 463
rect 446 468 450 472
rect 470 468 474 472
rect 486 468 490 472
rect 566 468 570 472
rect 734 468 738 472
rect 838 468 842 472
rect 846 468 850 472
rect 942 468 946 472
rect 982 468 986 472
rect 1078 468 1082 472
rect 1110 468 1114 472
rect 1174 468 1178 472
rect 1222 468 1226 472
rect 1246 468 1250 472
rect 1270 468 1274 472
rect 1350 468 1354 472
rect 1374 468 1378 472
rect 1398 468 1402 472
rect 1470 468 1474 472
rect 230 458 234 462
rect 270 458 274 462
rect 342 458 346 462
rect 374 458 378 462
rect 398 458 402 462
rect 406 458 410 462
rect 422 458 426 462
rect 462 458 466 462
rect 494 458 498 462
rect 598 459 602 463
rect 630 458 634 462
rect 670 458 674 462
rect 758 458 762 462
rect 782 458 786 462
rect 830 458 834 462
rect 862 458 866 462
rect 878 458 882 462
rect 886 458 890 462
rect 902 458 906 462
rect 910 458 914 462
rect 958 458 962 462
rect 966 458 970 462
rect 974 458 978 462
rect 1054 458 1058 462
rect 1070 458 1074 462
rect 1118 458 1122 462
rect 1126 458 1130 462
rect 1150 458 1154 462
rect 1182 458 1186 462
rect 1198 458 1202 462
rect 1238 458 1242 462
rect 1278 458 1282 462
rect 1286 458 1290 462
rect 1318 458 1322 462
rect 1358 458 1362 462
rect 1398 458 1402 462
rect 1430 458 1434 462
rect 1486 458 1490 462
rect 22 448 26 452
rect 86 448 90 452
rect 422 448 426 452
rect 782 448 786 452
rect 814 448 818 452
rect 1102 448 1106 452
rect 1142 448 1146 452
rect 1190 448 1194 452
rect 1294 448 1298 452
rect 1326 448 1330 452
rect 1414 448 1418 452
rect 62 438 66 442
rect 758 438 762 442
rect 1206 438 1210 442
rect 1310 438 1314 442
rect 1438 438 1442 442
rect 1478 438 1482 442
rect 926 418 930 422
rect 998 418 1002 422
rect 1086 418 1090 422
rect 1198 418 1202 422
rect 1262 418 1266 422
rect 1302 418 1306 422
rect 1318 418 1322 422
rect 1430 418 1434 422
rect 1502 418 1506 422
rect 490 403 494 407
rect 497 403 501 407
rect 278 388 282 392
rect 382 388 386 392
rect 462 388 466 392
rect 526 388 530 392
rect 638 388 642 392
rect 798 388 802 392
rect 1110 368 1114 372
rect 1286 368 1290 372
rect 1382 368 1386 372
rect 1454 368 1458 372
rect 70 358 74 362
rect 102 358 106 362
rect 166 358 170 362
rect 430 358 434 362
rect 454 358 458 362
rect 830 358 834 362
rect 862 358 866 362
rect 894 358 898 362
rect 982 358 986 362
rect 998 358 1002 362
rect 1094 358 1098 362
rect 1150 358 1154 362
rect 1190 358 1194 362
rect 1238 358 1242 362
rect 1302 358 1306 362
rect 1310 358 1314 362
rect 1390 358 1394 362
rect 1438 358 1442 362
rect 1470 358 1474 362
rect 38 348 42 352
rect 54 348 58 352
rect 118 348 122 352
rect 6 338 10 342
rect 62 338 66 342
rect 126 338 130 342
rect 214 347 218 351
rect 310 347 314 351
rect 374 348 378 352
rect 582 348 586 352
rect 670 347 674 351
rect 766 348 770 352
rect 814 348 818 352
rect 838 348 842 352
rect 878 348 882 352
rect 910 348 914 352
rect 918 348 922 352
rect 934 348 938 352
rect 974 348 978 352
rect 1046 348 1050 352
rect 1086 348 1090 352
rect 1102 348 1106 352
rect 1126 348 1130 352
rect 1134 348 1138 352
rect 1190 348 1194 352
rect 1222 348 1226 352
rect 1286 348 1290 352
rect 1318 348 1322 352
rect 1334 348 1338 352
rect 1366 348 1370 352
rect 1390 348 1394 352
rect 1406 348 1410 352
rect 182 338 186 342
rect 398 338 402 342
rect 446 338 450 342
rect 470 338 474 342
rect 486 338 490 342
rect 542 338 546 342
rect 94 328 98 332
rect 214 328 218 332
rect 310 328 314 332
rect 654 338 658 342
rect 742 338 746 342
rect 806 338 810 342
rect 886 338 890 342
rect 1446 348 1450 352
rect 1486 348 1490 352
rect 974 338 978 342
rect 1022 338 1026 342
rect 1038 338 1042 342
rect 1078 338 1082 342
rect 1126 338 1130 342
rect 1182 338 1186 342
rect 1206 338 1210 342
rect 1214 338 1218 342
rect 1246 338 1250 342
rect 1262 338 1266 342
rect 1342 338 1346 342
rect 1358 338 1362 342
rect 1414 338 1418 342
rect 1430 338 1434 342
rect 1502 338 1506 342
rect 574 328 578 332
rect 606 328 610 332
rect 766 328 770 332
rect 782 328 786 332
rect 790 328 794 332
rect 854 328 858 332
rect 894 328 898 332
rect 934 328 938 332
rect 1046 328 1050 332
rect 1070 328 1074 332
rect 1246 328 1250 332
rect 1390 328 1394 332
rect 1430 328 1434 332
rect 102 318 106 322
rect 734 318 738 322
rect 830 318 834 322
rect 846 318 850 322
rect 862 318 866 322
rect 958 318 962 322
rect 1166 318 1170 322
rect 1190 318 1194 322
rect 1254 318 1258 322
rect 1454 318 1458 322
rect 1470 318 1474 322
rect 1002 303 1006 307
rect 1009 303 1013 307
rect 222 288 226 292
rect 318 288 322 292
rect 414 288 418 292
rect 510 288 514 292
rect 622 288 626 292
rect 910 288 914 292
rect 1038 288 1042 292
rect 1470 288 1474 292
rect 838 278 842 282
rect 846 278 850 282
rect 854 278 858 282
rect 6 268 10 272
rect 78 268 82 272
rect 142 268 146 272
rect 238 268 242 272
rect 334 268 338 272
rect 574 268 578 272
rect 702 268 706 272
rect 774 268 778 272
rect 862 268 866 272
rect 902 278 906 282
rect 950 278 954 282
rect 1030 278 1034 282
rect 1102 278 1106 282
rect 1110 278 1114 282
rect 1134 278 1138 282
rect 1214 278 1218 282
rect 1262 278 1266 282
rect 1342 278 1346 282
rect 958 268 962 272
rect 974 268 978 272
rect 1046 268 1050 272
rect 1142 268 1146 272
rect 1166 268 1170 272
rect 1190 268 1194 272
rect 1206 268 1210 272
rect 1294 268 1298 272
rect 1310 268 1314 272
rect 1382 268 1386 272
rect 1430 268 1434 272
rect 1494 268 1498 272
rect 94 258 98 262
rect 158 259 162 263
rect 254 259 258 263
rect 350 259 354 263
rect 446 259 450 263
rect 478 258 482 262
rect 558 259 562 263
rect 870 258 874 262
rect 878 258 882 262
rect 926 258 930 262
rect 934 258 938 262
rect 974 258 978 262
rect 998 258 1002 262
rect 1054 258 1058 262
rect 1078 258 1082 262
rect 1086 258 1090 262
rect 1102 258 1106 262
rect 1126 258 1130 262
rect 1230 258 1234 262
rect 1262 258 1266 262
rect 1278 258 1282 262
rect 1318 258 1322 262
rect 1326 258 1330 262
rect 1342 258 1346 262
rect 1366 258 1370 262
rect 1390 258 1394 262
rect 1398 258 1402 262
rect 1446 258 1450 262
rect 1486 258 1490 262
rect 918 248 922 252
rect 1006 248 1010 252
rect 1254 248 1258 252
rect 1310 248 1314 252
rect 1374 248 1378 252
rect 1406 248 1410 252
rect 1414 248 1418 252
rect 1438 248 1442 252
rect 1470 248 1474 252
rect 206 238 210 242
rect 990 238 994 242
rect 1070 238 1074 242
rect 1358 238 1362 242
rect 1366 238 1370 242
rect 1454 238 1458 242
rect 998 228 1002 232
rect 1446 228 1450 232
rect 62 218 66 222
rect 638 218 642 222
rect 758 218 762 222
rect 798 218 802 222
rect 1062 218 1066 222
rect 1158 218 1162 222
rect 1422 218 1426 222
rect 490 203 494 207
rect 497 203 501 207
rect 94 188 98 192
rect 262 188 266 192
rect 302 188 306 192
rect 702 188 706 192
rect 1046 188 1050 192
rect 1286 188 1290 192
rect 1478 188 1482 192
rect 414 168 418 172
rect 606 168 610 172
rect 726 168 730 172
rect 958 168 962 172
rect 1038 168 1042 172
rect 1094 168 1098 172
rect 1262 168 1266 172
rect 1326 168 1330 172
rect 422 158 426 162
rect 766 158 770 162
rect 798 158 802 162
rect 942 158 946 162
rect 1022 158 1026 162
rect 1054 158 1058 162
rect 1078 158 1082 162
rect 1262 158 1266 162
rect 1494 158 1498 162
rect 54 148 58 152
rect 62 148 66 152
rect 198 147 202 151
rect 366 148 370 152
rect 438 148 442 152
rect 454 148 458 152
rect 478 148 482 152
rect 494 148 498 152
rect 542 147 546 151
rect 574 148 578 152
rect 646 148 650 152
rect 782 148 786 152
rect 822 148 826 152
rect 846 148 850 152
rect 934 148 938 152
rect 950 148 954 152
rect 974 148 978 152
rect 1046 148 1050 152
rect 1062 148 1066 152
rect 1094 148 1098 152
rect 1118 148 1122 152
rect 1166 148 1170 152
rect 1230 148 1234 152
rect 1254 148 1258 152
rect 1270 148 1274 152
rect 166 138 170 142
rect 206 138 210 142
rect 270 138 274 142
rect 318 138 322 142
rect 334 138 338 142
rect 454 138 458 142
rect 638 138 642 142
rect 710 138 714 142
rect 734 138 738 142
rect 774 138 778 142
rect 854 138 858 142
rect 878 140 882 144
rect 926 138 930 142
rect 1374 147 1378 151
rect 1470 148 1474 152
rect 1102 138 1106 142
rect 1110 138 1114 142
rect 1150 138 1154 142
rect 1222 138 1226 142
rect 1342 138 1346 142
rect 1358 138 1362 142
rect 1462 138 1466 142
rect 1470 138 1474 142
rect 102 128 106 132
rect 470 128 474 132
rect 542 128 546 132
rect 750 128 754 132
rect 822 128 826 132
rect 902 128 906 132
rect 918 128 922 132
rect 974 128 978 132
rect 1022 128 1026 132
rect 1070 128 1074 132
rect 1142 128 1146 132
rect 1206 128 1210 132
rect 1214 128 1218 132
rect 1238 128 1242 132
rect 110 118 114 122
rect 134 118 138 122
rect 798 118 802 122
rect 830 118 834 122
rect 862 118 866 122
rect 982 118 986 122
rect 1134 118 1138 122
rect 1246 118 1250 122
rect 1002 103 1006 107
rect 1009 103 1013 107
rect 38 88 42 92
rect 86 88 90 92
rect 150 88 154 92
rect 254 88 258 92
rect 318 88 322 92
rect 366 88 370 92
rect 510 88 514 92
rect 606 88 610 92
rect 1470 88 1474 92
rect 6 68 10 72
rect 54 68 58 72
rect 62 68 66 72
rect 110 68 114 72
rect 118 68 122 72
rect 166 68 170 72
rect 326 78 330 82
rect 342 78 346 82
rect 542 78 546 82
rect 910 78 914 82
rect 222 68 226 72
rect 270 68 274 72
rect 278 68 282 72
rect 302 68 306 72
rect 326 68 330 72
rect 350 68 354 72
rect 398 68 402 72
rect 446 68 450 72
rect 718 68 722 72
rect 806 68 810 72
rect 998 68 1002 72
rect 1118 68 1122 72
rect 1238 68 1242 72
rect 1358 68 1362 72
rect 1486 68 1490 72
rect 102 58 106 62
rect 190 58 194 62
rect 310 58 314 62
rect 430 59 434 63
rect 542 59 546 63
rect 550 58 554 62
rect 702 59 706 63
rect 822 59 826 63
rect 878 59 882 63
rect 62 48 66 52
rect 78 48 82 52
rect 86 48 90 52
rect 174 48 178 52
rect 1014 59 1018 63
rect 1134 59 1138 63
rect 1254 59 1258 63
rect 1382 58 1386 62
rect 1470 48 1474 52
rect 614 18 618 22
rect 734 18 738 22
rect 966 18 970 22
rect 1102 18 1106 22
rect 1222 18 1226 22
rect 1342 18 1346 22
rect 1462 18 1466 22
rect 490 3 494 7
rect 497 3 501 7
<< metal2 >>
rect 214 1328 218 1332
rect 238 1328 242 1332
rect 454 1328 458 1332
rect 478 1331 482 1332
rect 470 1328 482 1331
rect 10 1278 14 1281
rect 58 1278 62 1281
rect 22 1262 25 1268
rect 62 1262 65 1268
rect 78 1262 81 1278
rect 106 1268 110 1271
rect 86 1262 89 1268
rect 166 1262 169 1268
rect 74 1258 78 1261
rect 106 1258 110 1261
rect 138 1258 142 1261
rect 6 1252 9 1258
rect 38 1252 41 1258
rect 22 1162 25 1168
rect 6 1142 9 1148
rect 22 1142 25 1158
rect 78 1142 81 1148
rect 94 1142 97 1258
rect 174 1252 177 1288
rect 214 1282 217 1328
rect 238 1302 241 1328
rect 230 1298 238 1301
rect 230 1282 233 1298
rect 238 1272 241 1278
rect 286 1272 289 1298
rect 298 1288 302 1291
rect 202 1268 206 1271
rect 214 1262 217 1268
rect 310 1252 313 1268
rect 342 1263 345 1268
rect 266 1248 270 1251
rect 290 1248 294 1251
rect 170 1158 174 1161
rect 202 1158 206 1161
rect 266 1158 270 1161
rect 58 1118 62 1121
rect 14 1092 17 1108
rect 22 1102 25 1118
rect 70 1092 73 1118
rect 86 1112 89 1128
rect 102 1122 105 1148
rect 158 1142 161 1148
rect 178 1138 182 1141
rect 166 1122 169 1128
rect 38 1082 41 1088
rect 74 1078 78 1081
rect 6 1072 9 1078
rect 22 1072 25 1078
rect 22 1052 25 1058
rect 46 1052 49 1078
rect 86 1072 89 1098
rect 134 1063 137 1118
rect 190 1112 193 1148
rect 286 1142 289 1148
rect 210 1138 214 1141
rect 230 1132 233 1138
rect 202 1088 206 1091
rect 166 1062 169 1068
rect 102 1052 105 1058
rect 214 1052 217 1118
rect 294 1092 297 1098
rect 302 1072 305 1248
rect 318 1151 321 1158
rect 350 1152 353 1268
rect 374 1262 377 1268
rect 430 1262 433 1278
rect 454 1262 457 1328
rect 470 1282 473 1328
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1013 1303 1016 1307
rect 1070 1282 1073 1288
rect 482 1278 486 1281
rect 1474 1278 1478 1281
rect 470 1272 473 1278
rect 466 1258 470 1261
rect 414 1252 417 1258
rect 478 1252 481 1258
rect 438 1242 441 1248
rect 402 1218 406 1221
rect 394 1148 398 1151
rect 394 1128 398 1131
rect 406 1122 409 1128
rect 386 1118 390 1121
rect 422 1102 425 1218
rect 454 1192 457 1228
rect 430 1142 433 1148
rect 446 1142 449 1148
rect 442 1128 446 1131
rect 430 1122 433 1128
rect 410 1088 414 1091
rect 350 1072 353 1078
rect 358 1072 361 1088
rect 438 1082 441 1088
rect 462 1072 465 1238
rect 510 1232 513 1268
rect 526 1242 529 1248
rect 534 1232 537 1278
rect 614 1272 617 1278
rect 1062 1272 1065 1278
rect 1094 1272 1097 1278
rect 1174 1272 1177 1278
rect 810 1268 814 1271
rect 582 1242 585 1258
rect 598 1242 601 1268
rect 630 1252 633 1259
rect 488 1203 490 1207
rect 494 1203 497 1207
rect 501 1203 504 1207
rect 518 1162 521 1218
rect 530 1158 534 1161
rect 554 1158 558 1161
rect 542 1152 545 1158
rect 582 1152 585 1158
rect 482 1148 486 1151
rect 594 1148 598 1151
rect 654 1151 657 1158
rect 662 1142 665 1258
rect 694 1212 697 1218
rect 506 1138 510 1141
rect 546 1138 550 1141
rect 470 1132 473 1138
rect 558 1132 561 1138
rect 566 1132 569 1138
rect 618 1128 622 1131
rect 502 1072 505 1088
rect 362 1068 366 1071
rect 482 1068 486 1071
rect 230 1062 233 1068
rect 6 932 9 948
rect 22 942 25 948
rect 38 942 41 968
rect 94 962 97 1018
rect 134 952 137 958
rect 58 948 62 951
rect 198 951 201 958
rect 230 952 233 1058
rect 90 940 94 943
rect 30 932 33 938
rect 6 872 9 878
rect 50 868 54 871
rect 22 862 25 868
rect 38 852 41 868
rect 34 848 38 851
rect 22 842 25 848
rect 30 832 33 838
rect 70 832 73 928
rect 78 862 81 918
rect 110 892 113 918
rect 102 882 105 888
rect 118 882 121 938
rect 166 892 169 938
rect 138 878 142 881
rect 154 878 158 881
rect 186 878 190 881
rect 122 858 126 861
rect 78 842 81 848
rect 86 842 89 858
rect 106 848 110 851
rect 158 832 161 868
rect 174 852 177 868
rect 186 858 190 861
rect 6 732 9 778
rect 50 748 54 751
rect 38 742 41 748
rect 118 742 121 748
rect 22 732 25 738
rect 54 732 57 738
rect 94 732 98 735
rect 126 732 129 818
rect 174 762 177 848
rect 198 771 201 818
rect 190 768 201 771
rect 150 752 153 758
rect 138 748 142 751
rect 114 728 118 731
rect 6 682 9 728
rect 38 722 41 728
rect 18 718 22 721
rect 46 692 49 718
rect 22 672 25 678
rect 30 672 33 688
rect 94 682 97 718
rect 158 692 161 758
rect 182 742 185 758
rect 190 752 193 768
rect 206 742 209 938
rect 246 892 249 1058
rect 374 1052 377 1068
rect 430 1062 433 1068
rect 450 1058 454 1061
rect 466 1058 470 1061
rect 362 1048 366 1051
rect 450 1048 454 1051
rect 262 952 265 968
rect 278 942 281 1038
rect 302 942 305 948
rect 214 872 217 888
rect 310 882 313 938
rect 214 862 217 868
rect 278 852 281 868
rect 310 842 313 859
rect 226 747 230 750
rect 166 732 169 738
rect 206 732 209 738
rect 174 702 177 718
rect 214 692 217 708
rect 270 692 273 838
rect 286 762 289 768
rect 318 751 321 968
rect 326 692 329 1018
rect 374 1002 377 1048
rect 534 1042 537 1058
rect 488 1003 490 1007
rect 494 1003 497 1007
rect 501 1003 504 1007
rect 358 992 361 998
rect 542 992 545 1038
rect 550 981 553 1068
rect 566 1042 569 1128
rect 582 1052 585 1059
rect 542 978 553 981
rect 406 952 409 958
rect 386 948 390 951
rect 438 951 441 958
rect 466 948 470 951
rect 382 932 385 938
rect 406 932 409 938
rect 370 928 374 931
rect 370 918 374 921
rect 382 891 385 928
rect 526 922 529 928
rect 502 912 505 918
rect 378 888 385 891
rect 502 872 505 878
rect 406 863 409 868
rect 430 862 433 868
rect 482 858 486 861
rect 346 748 350 751
rect 126 682 129 688
rect 46 675 50 678
rect 130 678 137 681
rect 86 672 89 678
rect 106 668 110 671
rect 134 662 137 678
rect 150 662 153 678
rect 174 672 177 678
rect 286 672 289 678
rect 158 662 161 668
rect 18 658 22 661
rect 230 652 233 668
rect 238 662 241 668
rect 154 648 158 651
rect 294 642 297 668
rect 314 658 318 661
rect 38 552 41 558
rect 54 542 57 618
rect 126 592 129 618
rect 190 592 193 638
rect 314 588 318 591
rect 86 551 89 558
rect 86 492 89 528
rect 6 472 9 478
rect 46 475 50 478
rect 110 472 113 588
rect 246 562 249 568
rect 350 562 353 678
rect 238 552 241 558
rect 294 552 297 558
rect 266 548 270 551
rect 118 522 121 548
rect 326 542 329 548
rect 150 522 153 528
rect 166 472 169 478
rect 182 472 185 518
rect 22 452 25 468
rect 98 458 102 461
rect 138 458 142 461
rect 30 452 33 458
rect 62 442 65 458
rect 198 452 201 459
rect 82 448 86 451
rect 70 362 73 368
rect 98 358 102 361
rect 162 358 166 361
rect 6 342 9 358
rect 34 348 38 351
rect 54 342 57 348
rect 62 342 65 358
rect 182 352 185 418
rect 206 392 209 538
rect 214 532 217 538
rect 250 528 254 531
rect 262 492 265 528
rect 334 472 337 528
rect 358 482 361 708
rect 366 662 369 788
rect 414 751 417 758
rect 430 752 433 858
rect 518 852 521 859
rect 488 803 490 807
rect 494 803 497 807
rect 501 803 504 807
rect 430 742 433 748
rect 526 742 529 747
rect 378 738 382 741
rect 398 663 401 688
rect 430 672 433 738
rect 482 718 486 721
rect 494 672 497 678
rect 526 672 529 728
rect 430 662 433 668
rect 398 542 401 548
rect 422 542 425 548
rect 430 542 433 658
rect 510 652 513 659
rect 382 532 385 538
rect 462 522 465 618
rect 478 592 481 628
rect 488 603 490 607
rect 494 603 497 607
rect 501 603 504 607
rect 526 592 529 608
rect 542 582 545 978
rect 606 972 609 1128
rect 662 1072 665 1138
rect 662 1062 665 1068
rect 614 1052 617 1058
rect 650 1018 654 1021
rect 606 962 609 968
rect 582 942 585 958
rect 566 932 569 938
rect 590 932 593 948
rect 554 928 558 931
rect 598 931 601 958
rect 662 952 665 1038
rect 606 942 609 948
rect 634 938 638 941
rect 646 932 649 938
rect 594 928 601 931
rect 634 928 638 931
rect 566 821 569 928
rect 558 818 569 821
rect 574 882 577 918
rect 586 878 590 881
rect 550 592 553 618
rect 558 592 561 818
rect 574 792 577 878
rect 614 862 617 918
rect 630 892 633 918
rect 638 822 641 868
rect 586 818 590 821
rect 574 692 577 778
rect 638 772 641 778
rect 646 772 649 928
rect 662 902 665 948
rect 670 892 673 1018
rect 678 992 681 1148
rect 686 1052 689 1058
rect 702 1022 705 1268
rect 758 1242 761 1268
rect 790 1252 793 1258
rect 862 1242 865 1258
rect 730 1228 734 1231
rect 758 1192 761 1238
rect 790 1192 793 1218
rect 878 1202 881 1268
rect 934 1262 937 1268
rect 922 1258 926 1261
rect 886 1252 889 1258
rect 894 1231 897 1258
rect 902 1242 905 1258
rect 918 1242 921 1248
rect 894 1228 905 1231
rect 902 1192 905 1228
rect 942 1222 945 1268
rect 970 1258 977 1261
rect 958 1232 961 1238
rect 966 1222 969 1228
rect 910 1172 913 1218
rect 898 1168 902 1171
rect 814 1142 817 1158
rect 862 1152 865 1168
rect 902 1162 905 1168
rect 874 1158 878 1161
rect 882 1158 889 1161
rect 854 1142 857 1148
rect 794 1138 801 1141
rect 722 1118 726 1121
rect 750 1072 753 1132
rect 782 1092 785 1108
rect 798 1072 801 1138
rect 814 1092 817 1138
rect 810 1068 814 1071
rect 750 1042 753 1068
rect 798 1062 801 1068
rect 742 982 745 1018
rect 754 958 758 961
rect 706 948 710 951
rect 678 932 681 948
rect 686 942 689 948
rect 698 938 702 941
rect 718 932 721 958
rect 726 942 729 948
rect 678 892 681 928
rect 718 912 721 918
rect 734 911 737 948
rect 750 942 753 948
rect 766 932 769 958
rect 762 928 766 931
rect 774 921 777 1058
rect 822 1052 825 1118
rect 846 1092 849 1138
rect 886 1132 889 1158
rect 878 1082 881 1118
rect 894 1112 897 1158
rect 902 1142 905 1148
rect 902 1092 905 1138
rect 926 1132 929 1198
rect 942 1192 945 1218
rect 974 1212 977 1258
rect 982 1252 985 1268
rect 958 1192 961 1208
rect 982 1202 985 1248
rect 1006 1192 1009 1268
rect 934 1182 937 1188
rect 950 1172 953 1178
rect 958 1152 961 1158
rect 966 1142 969 1158
rect 990 1142 993 1158
rect 978 1138 982 1141
rect 998 1132 1001 1148
rect 926 1092 929 1128
rect 934 1092 937 1118
rect 974 1112 977 1128
rect 1014 1122 1017 1258
rect 1046 1192 1049 1258
rect 1046 1132 1049 1178
rect 1062 1132 1065 1238
rect 1070 1192 1073 1258
rect 1070 1152 1073 1188
rect 1078 1142 1081 1268
rect 1126 1262 1129 1268
rect 1098 1258 1102 1261
rect 1110 1212 1113 1258
rect 1118 1252 1121 1258
rect 1126 1182 1129 1188
rect 1142 1162 1145 1218
rect 1182 1172 1185 1258
rect 1190 1182 1193 1268
rect 1206 1162 1209 1278
rect 1214 1272 1217 1278
rect 1218 1258 1222 1261
rect 1230 1192 1233 1248
rect 1238 1232 1241 1258
rect 1262 1252 1265 1268
rect 1310 1242 1313 1268
rect 1350 1262 1353 1278
rect 1358 1272 1361 1278
rect 1378 1268 1382 1271
rect 1318 1252 1321 1258
rect 1250 1238 1254 1241
rect 1282 1238 1286 1241
rect 1326 1222 1329 1258
rect 1254 1192 1257 1218
rect 1334 1212 1337 1238
rect 1346 1228 1350 1231
rect 1366 1212 1369 1268
rect 1374 1222 1377 1258
rect 1390 1252 1393 1258
rect 1222 1172 1225 1178
rect 1246 1172 1249 1178
rect 1214 1152 1217 1168
rect 1262 1162 1265 1168
rect 1126 1142 1129 1148
rect 1242 1138 1246 1141
rect 1070 1122 1073 1138
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1013 1103 1016 1107
rect 922 1078 926 1081
rect 974 1078 982 1081
rect 838 1062 841 1068
rect 822 1022 825 1048
rect 830 1012 833 1058
rect 838 982 841 1058
rect 854 1042 857 1078
rect 874 1058 878 1061
rect 890 1048 894 1051
rect 890 1038 897 1041
rect 882 1028 886 1031
rect 870 992 873 998
rect 894 992 897 1038
rect 910 1041 913 1058
rect 918 1052 921 1078
rect 910 1038 921 1041
rect 902 1032 905 1038
rect 918 992 921 1038
rect 942 1032 945 1068
rect 950 1062 953 1068
rect 958 1052 961 1058
rect 966 1052 969 1068
rect 966 1022 969 1048
rect 974 1042 977 1078
rect 982 1062 985 1068
rect 990 1062 993 1068
rect 974 992 977 1038
rect 850 988 854 991
rect 998 982 1001 1018
rect 1014 992 1017 1088
rect 1150 1082 1153 1138
rect 1182 1122 1185 1135
rect 1198 1132 1201 1138
rect 1254 1132 1257 1148
rect 1278 1142 1281 1178
rect 1350 1152 1353 1198
rect 1358 1172 1361 1178
rect 1366 1172 1369 1208
rect 1374 1152 1377 1218
rect 1382 1162 1385 1238
rect 1398 1222 1401 1258
rect 1386 1158 1390 1161
rect 1386 1148 1390 1151
rect 1350 1142 1353 1148
rect 1398 1142 1401 1208
rect 1414 1202 1417 1268
rect 1438 1172 1441 1178
rect 1426 1168 1430 1171
rect 1290 1128 1294 1131
rect 1070 1062 1073 1068
rect 1094 1062 1097 1078
rect 1130 1068 1134 1071
rect 1154 1058 1161 1061
rect 1186 1058 1190 1061
rect 1202 1058 1206 1061
rect 1046 1052 1049 1058
rect 1078 1052 1081 1058
rect 794 968 798 971
rect 930 968 934 971
rect 854 962 857 968
rect 826 958 830 961
rect 726 908 737 911
rect 766 918 777 921
rect 834 948 838 951
rect 686 892 689 898
rect 726 892 729 908
rect 766 892 769 918
rect 654 882 657 888
rect 658 868 662 871
rect 678 852 681 868
rect 718 862 721 868
rect 710 852 713 858
rect 586 768 590 771
rect 602 768 606 771
rect 626 768 630 771
rect 618 758 622 761
rect 590 738 598 741
rect 590 722 593 738
rect 630 732 633 768
rect 646 752 649 758
rect 638 742 641 748
rect 662 742 665 848
rect 678 762 681 848
rect 686 842 689 848
rect 686 772 689 838
rect 674 748 678 751
rect 666 738 670 741
rect 638 721 641 738
rect 650 728 654 731
rect 630 718 641 721
rect 590 712 593 718
rect 582 602 585 668
rect 430 482 433 488
rect 438 482 441 518
rect 478 492 481 578
rect 590 572 593 708
rect 598 692 601 718
rect 606 672 609 688
rect 622 662 625 668
rect 618 648 622 651
rect 502 552 505 568
rect 558 562 561 568
rect 606 562 609 648
rect 630 572 633 718
rect 662 682 665 718
rect 682 678 689 681
rect 686 672 689 678
rect 646 662 649 668
rect 678 662 681 668
rect 694 662 697 678
rect 654 652 657 658
rect 638 622 641 638
rect 646 632 649 648
rect 670 622 673 638
rect 702 632 705 758
rect 710 752 713 848
rect 734 842 737 868
rect 742 831 745 858
rect 734 828 745 831
rect 718 752 721 758
rect 726 742 729 768
rect 734 752 737 828
rect 758 792 761 888
rect 774 862 777 868
rect 766 842 769 848
rect 790 772 793 848
rect 798 762 801 948
rect 834 938 838 941
rect 806 892 809 938
rect 838 872 841 878
rect 810 868 814 871
rect 826 868 830 871
rect 822 852 825 858
rect 838 762 841 868
rect 846 862 849 918
rect 862 912 865 938
rect 862 892 865 898
rect 870 882 873 968
rect 942 962 945 968
rect 958 962 961 978
rect 890 958 894 961
rect 962 958 966 961
rect 986 958 990 961
rect 878 952 881 958
rect 1014 952 1017 968
rect 902 922 905 938
rect 918 922 921 948
rect 902 882 905 908
rect 918 892 921 918
rect 846 782 849 858
rect 854 762 857 768
rect 746 748 750 751
rect 770 748 774 751
rect 802 748 806 751
rect 702 592 705 598
rect 546 558 550 561
rect 586 558 590 561
rect 510 542 513 548
rect 526 532 529 558
rect 606 552 609 558
rect 546 548 550 551
rect 566 542 569 548
rect 614 542 617 568
rect 630 562 633 568
rect 586 538 590 541
rect 618 538 622 541
rect 534 492 537 538
rect 630 532 633 558
rect 638 552 641 558
rect 662 552 665 568
rect 710 551 713 728
rect 734 712 737 748
rect 734 672 737 678
rect 718 642 721 658
rect 718 562 721 638
rect 726 612 729 658
rect 742 572 745 748
rect 838 742 841 758
rect 854 752 857 758
rect 862 752 865 878
rect 914 868 918 871
rect 870 812 873 868
rect 894 852 897 858
rect 894 842 897 848
rect 886 822 889 828
rect 854 742 857 748
rect 862 742 865 748
rect 870 742 873 808
rect 918 762 921 768
rect 918 752 921 758
rect 934 752 937 948
rect 1010 938 1014 941
rect 942 932 945 938
rect 966 892 969 938
rect 966 882 969 888
rect 974 872 977 908
rect 990 872 993 938
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1013 903 1016 907
rect 946 868 950 871
rect 978 868 982 871
rect 958 862 961 868
rect 942 832 945 848
rect 950 812 953 858
rect 962 818 966 821
rect 958 752 961 758
rect 966 752 969 798
rect 930 748 934 751
rect 894 742 897 748
rect 918 742 921 748
rect 794 738 798 741
rect 706 548 713 551
rect 742 552 745 558
rect 638 522 641 548
rect 654 542 657 548
rect 686 542 689 548
rect 718 538 726 541
rect 746 538 750 541
rect 758 541 761 718
rect 774 672 777 678
rect 822 672 825 708
rect 794 668 798 671
rect 794 658 798 661
rect 766 652 769 658
rect 774 652 777 658
rect 810 648 814 651
rect 790 642 793 648
rect 802 638 806 641
rect 774 552 777 618
rect 798 572 801 628
rect 774 542 777 548
rect 822 542 825 668
rect 838 552 841 678
rect 846 552 849 698
rect 854 682 857 718
rect 870 692 873 738
rect 758 538 766 541
rect 582 512 585 518
rect 446 482 449 488
rect 606 482 609 518
rect 630 502 633 518
rect 346 478 350 481
rect 398 472 401 478
rect 230 462 233 468
rect 274 458 278 461
rect 274 388 278 391
rect 114 348 118 351
rect 214 351 217 358
rect 126 342 129 348
rect 182 342 185 348
rect 94 332 97 338
rect 102 278 105 318
rect 214 272 217 328
rect 222 292 225 388
rect 310 342 313 347
rect 310 272 313 328
rect 318 292 321 458
rect 334 442 337 468
rect 422 462 425 468
rect 346 458 350 461
rect 378 458 382 461
rect 394 458 398 461
rect 406 452 409 458
rect 426 448 430 451
rect 382 392 385 448
rect 426 358 430 361
rect 374 352 377 358
rect 446 342 449 468
rect 462 462 465 478
rect 566 472 569 478
rect 482 468 486 471
rect 470 462 473 468
rect 458 458 462 461
rect 490 458 494 461
rect 462 392 465 448
rect 598 432 601 459
rect 626 458 630 461
rect 646 432 649 518
rect 662 492 665 528
rect 694 502 697 538
rect 662 472 665 488
rect 694 462 697 498
rect 674 458 678 461
rect 702 442 705 448
rect 488 403 490 407
rect 494 403 497 407
rect 501 403 504 407
rect 526 392 529 428
rect 638 392 641 408
rect 454 362 457 368
rect 486 342 489 358
rect 670 351 673 358
rect 398 292 401 338
rect 410 288 414 291
rect 334 272 337 278
rect 10 268 14 271
rect 74 268 78 271
rect 38 92 41 268
rect 94 252 97 258
rect 142 242 145 268
rect 158 252 161 259
rect 206 242 209 268
rect 238 262 241 268
rect 62 222 65 238
rect 62 152 65 218
rect 54 72 57 148
rect 86 92 89 228
rect 94 192 97 218
rect 166 142 169 148
rect 198 142 201 147
rect 206 142 209 238
rect 106 128 110 131
rect 138 118 142 121
rect 66 68 70 71
rect 6 52 9 68
rect 102 62 105 78
rect 110 72 113 118
rect 118 72 121 118
rect 150 92 153 118
rect 166 82 169 138
rect 254 122 257 259
rect 262 192 265 238
rect 302 192 305 258
rect 334 142 337 268
rect 350 252 353 259
rect 446 222 449 259
rect 414 152 417 168
rect 422 162 425 168
rect 470 162 473 338
rect 542 332 545 338
rect 514 288 518 291
rect 478 262 481 268
rect 488 203 490 207
rect 494 203 497 207
rect 501 203 504 207
rect 494 152 497 158
rect 450 148 454 151
rect 482 148 486 151
rect 270 92 273 138
rect 318 92 321 138
rect 366 92 369 148
rect 438 142 441 148
rect 454 132 457 138
rect 466 128 470 131
rect 510 92 513 278
rect 574 272 577 328
rect 582 282 585 348
rect 606 332 609 338
rect 654 332 657 338
rect 626 288 630 291
rect 702 272 705 438
rect 574 262 577 268
rect 558 242 561 259
rect 574 152 577 258
rect 610 168 614 171
rect 542 142 545 147
rect 574 142 577 148
rect 250 88 254 91
rect 542 82 545 128
rect 606 92 609 148
rect 638 142 641 218
rect 698 188 702 191
rect 646 142 649 148
rect 330 78 334 81
rect 302 72 305 78
rect 166 62 169 68
rect 194 58 198 61
rect 78 52 81 58
rect 66 48 70 51
rect 86 42 89 48
rect 102 -18 105 58
rect 178 48 182 51
rect 102 -22 106 -18
rect 222 -19 225 68
rect 270 62 273 68
rect 278 52 281 68
rect 326 62 329 68
rect 342 62 345 78
rect 350 72 353 78
rect 446 72 449 78
rect 314 58 318 61
rect 238 -19 242 -18
rect 222 -22 242 -19
rect 350 -19 353 68
rect 398 62 401 68
rect 434 59 438 62
rect 550 62 553 68
rect 702 63 705 178
rect 710 142 713 308
rect 718 292 721 538
rect 802 528 806 531
rect 818 528 822 531
rect 838 522 841 538
rect 786 518 790 521
rect 726 342 729 518
rect 738 478 742 481
rect 758 471 761 518
rect 806 482 809 488
rect 814 482 817 488
rect 758 468 769 471
rect 734 452 737 468
rect 754 458 758 461
rect 754 438 758 441
rect 766 362 769 468
rect 778 458 782 461
rect 822 461 825 508
rect 830 502 833 518
rect 846 472 849 478
rect 822 458 830 461
rect 786 448 790 451
rect 810 448 814 451
rect 798 392 801 418
rect 738 338 742 341
rect 726 172 729 338
rect 738 318 742 321
rect 726 162 729 168
rect 734 142 737 148
rect 750 142 753 358
rect 806 352 809 358
rect 814 352 817 378
rect 766 342 769 348
rect 806 342 809 348
rect 778 328 782 331
rect 750 132 753 138
rect 718 72 721 78
rect 758 72 761 218
rect 766 182 769 328
rect 790 322 793 328
rect 774 272 777 278
rect 766 162 769 168
rect 798 162 801 218
rect 822 192 825 448
rect 838 432 841 468
rect 854 452 857 658
rect 870 542 873 548
rect 878 542 881 718
rect 886 652 889 738
rect 902 732 905 738
rect 914 728 918 731
rect 910 702 913 728
rect 934 682 937 688
rect 910 672 913 678
rect 942 672 945 718
rect 898 668 902 671
rect 918 662 921 668
rect 902 652 905 658
rect 934 652 937 658
rect 938 648 950 651
rect 886 632 889 648
rect 902 542 905 568
rect 910 552 913 588
rect 918 532 921 558
rect 926 552 929 588
rect 958 572 961 658
rect 966 622 969 748
rect 974 742 977 858
rect 982 762 985 858
rect 990 792 993 868
rect 1014 852 1017 868
rect 1022 862 1025 1048
rect 1034 1038 1038 1041
rect 1038 1022 1041 1038
rect 1046 1032 1049 1038
rect 1054 1012 1057 1048
rect 1086 1042 1089 1048
rect 1110 1042 1113 1048
rect 1066 1038 1070 1041
rect 1086 982 1089 1038
rect 1106 1028 1110 1031
rect 1118 992 1121 1048
rect 1150 1042 1153 1048
rect 1126 982 1129 1018
rect 1030 952 1033 978
rect 1090 968 1094 971
rect 1122 968 1126 971
rect 1030 892 1033 938
rect 1038 932 1041 938
rect 1038 912 1041 918
rect 998 782 1001 818
rect 1006 772 1009 848
rect 1014 752 1017 838
rect 990 732 993 738
rect 986 728 990 731
rect 1014 722 1017 748
rect 1022 742 1025 768
rect 1038 742 1041 908
rect 1046 892 1049 948
rect 1054 942 1057 958
rect 1074 948 1078 951
rect 1102 942 1105 958
rect 1066 938 1070 941
rect 1110 941 1113 958
rect 1118 952 1121 958
rect 1158 952 1161 1058
rect 1166 1032 1169 1048
rect 1178 1038 1182 1041
rect 1190 1032 1193 1048
rect 1198 1032 1201 1048
rect 1214 1042 1217 1068
rect 1230 1032 1233 1078
rect 1254 1072 1257 1128
rect 1302 1122 1305 1138
rect 1414 1132 1417 1158
rect 1438 1142 1441 1148
rect 1414 1122 1417 1128
rect 1286 1072 1289 1118
rect 1334 1082 1337 1118
rect 1342 1092 1345 1118
rect 1406 1092 1409 1118
rect 1282 1058 1286 1061
rect 1246 1032 1249 1058
rect 1294 1052 1297 1058
rect 1258 1048 1262 1051
rect 1274 1038 1278 1041
rect 1166 962 1169 1028
rect 1174 952 1177 1018
rect 1110 938 1121 941
rect 1066 928 1070 931
rect 1046 872 1049 888
rect 1110 882 1113 888
rect 1106 878 1110 881
rect 1054 842 1057 848
rect 1062 772 1065 858
rect 1070 852 1073 878
rect 1094 862 1097 868
rect 1110 862 1113 868
rect 1086 852 1089 858
rect 1118 852 1121 938
rect 1142 912 1145 948
rect 1150 942 1153 948
rect 1190 942 1193 968
rect 1230 962 1233 1028
rect 1238 972 1241 978
rect 1218 958 1222 961
rect 1218 948 1222 951
rect 1166 932 1169 938
rect 1190 932 1193 938
rect 1198 932 1201 948
rect 1230 932 1233 958
rect 1246 952 1249 1008
rect 1278 992 1281 998
rect 1270 972 1273 978
rect 1286 972 1289 1018
rect 1254 962 1257 968
rect 1242 948 1246 951
rect 1274 948 1278 951
rect 1126 862 1129 868
rect 1142 861 1145 908
rect 1166 872 1169 878
rect 1154 868 1158 871
rect 1142 858 1150 861
rect 1078 772 1081 818
rect 1110 762 1113 848
rect 1118 802 1121 848
rect 1134 832 1137 838
rect 1174 832 1177 878
rect 1182 852 1185 868
rect 1190 862 1193 928
rect 1206 892 1209 928
rect 1286 922 1289 958
rect 1294 922 1297 1048
rect 1302 1012 1305 1058
rect 1310 982 1313 1068
rect 1326 1062 1329 1078
rect 1366 1072 1369 1088
rect 1414 1072 1417 1078
rect 1422 1072 1425 1088
rect 1306 968 1310 971
rect 1318 962 1321 988
rect 1330 968 1334 971
rect 1342 962 1345 1028
rect 1350 1002 1353 1068
rect 1430 1062 1433 1068
rect 1446 1062 1449 1118
rect 1454 1082 1457 1188
rect 1462 1162 1465 1268
rect 1486 1162 1489 1218
rect 1462 1122 1465 1128
rect 1470 1122 1473 1128
rect 1358 992 1361 1058
rect 1382 1052 1385 1058
rect 1310 952 1313 958
rect 1366 952 1369 1048
rect 1374 972 1377 998
rect 1390 962 1393 988
rect 1406 972 1409 998
rect 1338 948 1342 951
rect 1394 948 1398 951
rect 1342 932 1345 938
rect 1218 878 1222 881
rect 1126 781 1129 818
rect 1182 792 1185 838
rect 1206 832 1209 858
rect 1206 782 1209 828
rect 1214 822 1217 868
rect 1238 862 1241 888
rect 1262 862 1265 868
rect 1270 862 1273 868
rect 1302 862 1305 918
rect 1318 892 1321 918
rect 1310 852 1313 878
rect 1322 868 1326 871
rect 1354 858 1358 861
rect 1238 842 1241 848
rect 1246 832 1249 848
rect 1302 842 1305 848
rect 1334 842 1337 858
rect 1366 852 1369 918
rect 1414 882 1417 918
rect 1422 892 1425 1048
rect 1438 972 1441 1058
rect 1446 1052 1449 1058
rect 1454 1041 1457 1078
rect 1478 1072 1481 1118
rect 1486 1102 1489 1138
rect 1494 1102 1497 1148
rect 1502 1092 1505 1258
rect 1494 1072 1497 1078
rect 1466 1058 1470 1061
rect 1474 1058 1486 1061
rect 1482 1048 1486 1051
rect 1454 1038 1462 1041
rect 1470 962 1473 1018
rect 1482 968 1486 971
rect 1502 962 1505 1068
rect 1510 1052 1513 1078
rect 1502 952 1505 958
rect 1490 948 1494 951
rect 1470 942 1473 948
rect 1458 938 1462 941
rect 1430 932 1433 938
rect 1430 892 1433 928
rect 1438 902 1441 918
rect 1446 882 1449 928
rect 1410 868 1414 871
rect 1430 862 1433 878
rect 1366 842 1369 848
rect 1382 842 1385 858
rect 1390 852 1393 858
rect 1438 852 1441 878
rect 1462 872 1465 918
rect 1478 862 1481 888
rect 1450 858 1454 861
rect 1466 848 1470 851
rect 1398 842 1401 848
rect 1486 842 1489 878
rect 1458 838 1462 841
rect 1350 832 1353 838
rect 1262 782 1265 818
rect 1126 778 1137 781
rect 1122 768 1126 771
rect 1134 762 1137 778
rect 1286 781 1289 818
rect 1302 792 1305 828
rect 1358 812 1361 818
rect 1390 802 1393 818
rect 1278 778 1289 781
rect 1390 782 1393 788
rect 1142 762 1145 778
rect 1154 768 1158 771
rect 1110 752 1113 758
rect 1134 752 1137 758
rect 1166 752 1169 758
rect 1082 748 1086 751
rect 1090 738 1094 741
rect 1070 732 1073 738
rect 1110 732 1113 748
rect 1126 742 1129 748
rect 1190 742 1193 778
rect 1278 772 1281 778
rect 1398 772 1401 778
rect 1414 772 1417 808
rect 1218 768 1222 771
rect 1198 732 1201 758
rect 1226 748 1230 751
rect 1206 742 1209 748
rect 1238 742 1241 768
rect 1286 762 1289 768
rect 1382 762 1385 768
rect 1314 758 1318 761
rect 1250 738 1254 741
rect 1262 732 1265 758
rect 1270 752 1273 758
rect 1290 738 1294 741
rect 1042 728 1046 731
rect 1058 728 1062 731
rect 1250 728 1254 731
rect 982 681 985 718
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1013 703 1016 707
rect 1030 692 1033 718
rect 974 678 985 681
rect 974 662 977 678
rect 990 671 993 688
rect 1078 682 1081 718
rect 1078 672 1081 678
rect 1110 672 1113 718
rect 1126 692 1129 728
rect 1130 678 1134 681
rect 986 668 993 671
rect 1030 652 1033 668
rect 1062 662 1065 668
rect 1150 662 1153 678
rect 1158 662 1161 718
rect 1198 692 1201 728
rect 1190 662 1193 678
rect 1206 672 1209 728
rect 1214 682 1217 718
rect 1266 688 1273 691
rect 1262 682 1265 688
rect 1246 672 1249 678
rect 1254 672 1257 678
rect 1042 658 1046 661
rect 1102 652 1105 658
rect 1206 652 1209 668
rect 1214 662 1217 668
rect 1034 648 1046 651
rect 1178 648 1182 651
rect 1194 648 1198 651
rect 1142 642 1145 648
rect 1158 642 1161 648
rect 1222 642 1225 668
rect 1234 658 1238 661
rect 1270 652 1273 688
rect 1282 658 1286 661
rect 1302 652 1305 748
rect 1310 662 1313 758
rect 1390 752 1393 768
rect 1410 758 1414 761
rect 1422 752 1425 768
rect 1298 648 1302 651
rect 1314 648 1318 651
rect 1286 642 1289 648
rect 938 568 942 571
rect 942 552 945 558
rect 958 552 961 568
rect 982 561 985 608
rect 990 572 993 618
rect 1062 592 1065 618
rect 1086 612 1089 618
rect 1086 588 1094 591
rect 1038 572 1041 578
rect 1066 568 1070 571
rect 1070 562 1073 568
rect 978 558 985 561
rect 1050 558 1054 561
rect 982 552 985 558
rect 966 532 969 548
rect 990 542 993 548
rect 1014 542 1017 548
rect 1026 538 1030 541
rect 882 528 886 531
rect 870 522 873 528
rect 898 518 902 521
rect 966 512 969 518
rect 870 492 873 508
rect 926 492 929 508
rect 866 478 870 481
rect 874 478 886 481
rect 942 472 945 478
rect 974 472 977 538
rect 1010 528 1014 531
rect 990 518 998 521
rect 982 492 985 498
rect 982 472 985 488
rect 990 482 993 518
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1013 503 1016 507
rect 1038 492 1041 528
rect 1054 522 1057 558
rect 1078 552 1081 578
rect 1086 562 1089 588
rect 1094 552 1097 588
rect 1102 542 1105 578
rect 1078 532 1081 538
rect 1118 532 1121 568
rect 1126 562 1129 588
rect 1150 582 1153 618
rect 1134 552 1137 578
rect 1146 568 1150 571
rect 1110 512 1113 518
rect 1030 482 1033 488
rect 1006 472 1009 478
rect 1070 472 1073 478
rect 1078 472 1081 488
rect 1110 472 1113 478
rect 862 462 865 468
rect 902 462 905 468
rect 974 462 977 468
rect 1070 462 1073 468
rect 1118 462 1121 498
rect 1142 482 1145 548
rect 1150 492 1153 518
rect 1166 492 1169 568
rect 1174 552 1177 618
rect 1310 592 1313 618
rect 1326 602 1329 738
rect 1374 732 1377 738
rect 1382 692 1385 748
rect 1430 692 1433 818
rect 1446 772 1449 818
rect 1458 768 1462 771
rect 1470 762 1473 838
rect 1486 832 1489 838
rect 1478 772 1481 818
rect 1494 762 1497 948
rect 1502 792 1505 938
rect 1510 902 1513 1048
rect 1458 748 1462 751
rect 1470 741 1473 758
rect 1478 752 1481 758
rect 1486 742 1489 748
rect 1470 738 1481 741
rect 1386 678 1390 681
rect 1338 658 1342 661
rect 1334 642 1337 648
rect 1350 642 1353 648
rect 1366 642 1369 658
rect 1374 652 1377 668
rect 1438 662 1441 718
rect 1418 658 1422 661
rect 1426 648 1430 651
rect 1438 642 1441 658
rect 1406 632 1409 638
rect 1298 578 1302 581
rect 1238 572 1241 578
rect 1182 562 1185 568
rect 1230 562 1233 568
rect 1246 562 1249 568
rect 1234 548 1238 551
rect 1190 542 1193 548
rect 1174 532 1177 538
rect 1198 532 1201 538
rect 1254 532 1257 558
rect 1278 552 1281 568
rect 1310 562 1313 568
rect 1282 548 1286 551
rect 1270 542 1273 548
rect 1294 542 1297 548
rect 1286 532 1289 538
rect 1218 528 1222 531
rect 1154 478 1158 481
rect 890 458 894 461
rect 830 332 833 358
rect 838 352 841 378
rect 862 352 865 358
rect 878 352 881 458
rect 890 358 894 361
rect 902 351 905 458
rect 910 452 913 458
rect 958 452 961 458
rect 910 352 913 358
rect 926 352 929 418
rect 934 352 937 448
rect 902 348 910 351
rect 854 332 857 348
rect 878 342 881 348
rect 918 342 921 348
rect 890 338 894 341
rect 830 272 833 318
rect 846 282 849 318
rect 862 302 865 318
rect 870 281 873 328
rect 862 278 873 281
rect 838 262 841 278
rect 854 272 857 278
rect 862 272 865 278
rect 870 262 873 268
rect 878 262 881 338
rect 934 332 937 338
rect 894 322 897 328
rect 910 292 913 328
rect 902 282 905 288
rect 934 262 937 318
rect 958 312 961 318
rect 946 278 950 281
rect 954 268 958 271
rect 966 261 969 458
rect 1054 452 1057 458
rect 1102 452 1105 458
rect 998 362 1001 418
rect 974 352 977 358
rect 974 332 977 338
rect 982 271 985 358
rect 1038 342 1041 448
rect 1086 361 1089 418
rect 1086 358 1094 361
rect 1086 352 1089 358
rect 1050 348 1054 351
rect 1098 348 1102 351
rect 1110 342 1113 368
rect 1126 362 1129 458
rect 1142 452 1145 478
rect 1170 468 1174 471
rect 1150 462 1153 468
rect 1198 462 1201 518
rect 1206 481 1209 518
rect 1230 492 1233 528
rect 1262 522 1265 528
rect 1206 478 1217 481
rect 1178 458 1182 461
rect 1190 452 1193 458
rect 1206 442 1209 468
rect 1134 352 1137 368
rect 1186 358 1190 361
rect 1150 352 1153 358
rect 1122 348 1126 351
rect 1026 338 1030 341
rect 1074 338 1078 341
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1013 303 1016 307
rect 1034 288 1038 291
rect 1046 282 1049 328
rect 1070 322 1073 328
rect 1102 282 1105 308
rect 1110 282 1113 288
rect 978 268 985 271
rect 966 258 974 261
rect 914 248 918 251
rect 926 172 929 258
rect 982 241 985 268
rect 994 258 998 261
rect 1006 252 1009 278
rect 1030 272 1033 278
rect 1118 272 1121 348
rect 1126 332 1129 338
rect 1134 312 1137 348
rect 1182 342 1185 358
rect 1198 351 1201 418
rect 1194 348 1201 351
rect 1198 341 1201 348
rect 1214 342 1217 478
rect 1222 442 1225 468
rect 1238 462 1241 488
rect 1250 468 1254 471
rect 1262 442 1265 478
rect 1270 472 1273 508
rect 1278 462 1281 528
rect 1242 358 1246 361
rect 1262 352 1265 418
rect 1286 372 1289 458
rect 1294 452 1297 538
rect 1310 472 1313 558
rect 1334 552 1337 628
rect 1342 552 1345 618
rect 1398 611 1401 618
rect 1390 608 1401 611
rect 1350 562 1353 568
rect 1358 552 1361 578
rect 1370 568 1374 571
rect 1334 541 1337 548
rect 1334 538 1345 541
rect 1322 518 1326 521
rect 1310 442 1313 468
rect 1318 462 1321 488
rect 1334 482 1337 508
rect 1342 492 1345 538
rect 1382 532 1385 538
rect 1374 492 1377 518
rect 1350 472 1353 488
rect 1366 462 1369 478
rect 1378 468 1382 471
rect 1326 442 1329 448
rect 1358 442 1361 458
rect 1302 362 1305 418
rect 1226 348 1230 351
rect 1198 338 1206 341
rect 1130 278 1134 281
rect 1046 252 1049 268
rect 1078 262 1081 268
rect 1126 262 1129 278
rect 1142 272 1145 298
rect 1166 292 1169 318
rect 1058 258 1062 261
rect 1090 258 1094 261
rect 982 238 990 241
rect 998 232 1001 248
rect 1070 242 1073 248
rect 1046 182 1049 188
rect 954 168 958 171
rect 1034 168 1038 171
rect 778 148 782 151
rect 842 148 846 151
rect 822 142 825 148
rect 854 142 857 158
rect 770 138 774 141
rect 926 142 929 168
rect 1022 162 1025 168
rect 1054 162 1057 198
rect 1062 162 1065 218
rect 1094 172 1097 178
rect 934 152 937 158
rect 942 152 945 158
rect 950 152 953 158
rect 1050 148 1054 151
rect 1058 148 1062 151
rect 974 142 977 148
rect 854 132 857 138
rect 826 128 830 131
rect 798 122 801 128
rect 878 122 881 140
rect 902 132 905 138
rect 918 132 921 138
rect 1022 132 1025 138
rect 1070 132 1073 158
rect 1078 142 1081 158
rect 1094 152 1097 158
rect 1102 152 1105 258
rect 1102 142 1105 148
rect 1110 142 1113 188
rect 1118 152 1121 168
rect 1150 162 1153 288
rect 1190 282 1193 318
rect 1214 282 1217 338
rect 1170 268 1174 271
rect 1202 268 1206 271
rect 1190 242 1193 268
rect 1230 262 1233 348
rect 1242 338 1246 341
rect 1258 338 1262 341
rect 1158 202 1161 218
rect 1246 192 1249 328
rect 1254 322 1257 328
rect 1258 278 1262 281
rect 1254 252 1257 268
rect 1262 172 1265 258
rect 1150 142 1153 158
rect 1162 148 1166 151
rect 1222 142 1225 168
rect 1254 152 1257 158
rect 1234 148 1238 151
rect 1262 142 1265 158
rect 1270 152 1273 278
rect 1278 262 1281 348
rect 1286 272 1289 348
rect 1310 292 1313 358
rect 1318 352 1321 418
rect 1334 352 1337 358
rect 1294 272 1297 288
rect 1334 282 1337 348
rect 1358 342 1361 418
rect 1366 352 1369 358
rect 1342 332 1345 338
rect 1342 282 1345 328
rect 1314 268 1318 271
rect 1294 262 1297 268
rect 1366 262 1369 268
rect 1330 258 1334 261
rect 1310 252 1313 258
rect 1318 252 1321 258
rect 1286 192 1289 218
rect 1326 152 1329 168
rect 1342 142 1345 258
rect 1374 252 1377 458
rect 1382 372 1385 418
rect 1390 362 1393 608
rect 1398 562 1401 598
rect 1430 592 1433 618
rect 1446 582 1449 658
rect 1454 652 1457 718
rect 1478 692 1481 738
rect 1502 732 1505 738
rect 1462 672 1465 678
rect 1398 542 1401 548
rect 1470 542 1473 588
rect 1486 572 1489 578
rect 1494 561 1497 618
rect 1510 602 1513 668
rect 1494 558 1502 561
rect 1482 548 1486 551
rect 1410 538 1414 541
rect 1482 538 1486 541
rect 1406 471 1409 518
rect 1454 492 1457 518
rect 1402 468 1409 471
rect 1454 472 1457 478
rect 1470 472 1473 538
rect 1470 462 1473 468
rect 1486 462 1489 468
rect 1398 452 1401 458
rect 1414 452 1417 458
rect 1430 452 1433 458
rect 1442 438 1446 441
rect 1430 361 1433 418
rect 1458 368 1462 371
rect 1470 362 1473 438
rect 1430 358 1438 361
rect 1386 348 1390 351
rect 1442 348 1446 351
rect 1478 351 1481 438
rect 1478 348 1486 351
rect 1406 342 1409 348
rect 1430 342 1433 348
rect 1390 332 1393 338
rect 1414 322 1417 338
rect 1426 328 1430 331
rect 1434 268 1438 271
rect 1382 262 1385 268
rect 1446 262 1449 308
rect 1454 272 1457 318
rect 1470 312 1473 318
rect 1470 292 1473 298
rect 1354 238 1358 241
rect 1366 232 1369 238
rect 1390 222 1393 258
rect 1398 252 1401 258
rect 1434 248 1438 251
rect 1466 248 1470 251
rect 1406 232 1409 248
rect 1414 242 1417 248
rect 1446 232 1449 238
rect 1374 151 1377 158
rect 1142 132 1145 138
rect 1206 132 1209 138
rect 970 128 974 131
rect 1234 128 1238 131
rect 1214 122 1217 128
rect 830 101 833 118
rect 822 98 833 101
rect 802 68 806 71
rect 822 63 825 98
rect 430 -18 433 59
rect 488 3 490 7
rect 494 3 497 7
rect 501 3 504 7
rect 542 -18 545 59
rect 862 62 865 118
rect 910 72 913 78
rect 878 63 881 68
rect 982 62 985 118
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1013 103 1016 107
rect 998 72 1001 78
rect 1118 72 1121 78
rect 1014 63 1017 68
rect 1134 63 1137 118
rect 1246 101 1249 118
rect 1246 98 1257 101
rect 1238 72 1241 78
rect 1254 63 1257 98
rect 1358 82 1361 138
rect 1358 72 1361 78
rect 1422 62 1425 218
rect 1454 132 1457 238
rect 1478 201 1481 348
rect 1494 272 1497 548
rect 1502 342 1505 418
rect 1486 262 1489 268
rect 1470 198 1481 201
rect 1470 152 1473 198
rect 1478 182 1481 188
rect 1490 158 1494 161
rect 1462 142 1465 148
rect 1474 138 1478 141
rect 1470 92 1473 128
rect 1486 72 1489 158
rect 1502 142 1505 338
rect 1386 58 1390 61
rect 1470 52 1473 58
rect 358 -19 362 -18
rect 350 -22 362 -19
rect 430 -22 434 -18
rect 542 -22 546 -18
rect 614 -19 617 18
rect 622 -19 626 -18
rect 614 -22 626 -19
rect 734 -19 737 18
rect 742 -19 746 -18
rect 734 -22 746 -19
rect 958 -19 962 -18
rect 966 -19 969 18
rect 958 -22 969 -19
rect 1094 -19 1098 -18
rect 1102 -19 1105 18
rect 1094 -22 1105 -19
rect 1214 -19 1218 -18
rect 1222 -19 1225 18
rect 1214 -22 1225 -19
rect 1334 -19 1338 -18
rect 1342 -19 1345 18
rect 1334 -22 1345 -19
rect 1454 -19 1458 -18
rect 1462 -19 1465 18
rect 1454 -22 1465 -19
<< m3contact >>
rect 174 1288 178 1292
rect 14 1278 18 1282
rect 54 1278 58 1282
rect 22 1268 26 1272
rect 110 1268 114 1272
rect 166 1268 170 1272
rect 62 1258 66 1262
rect 70 1258 74 1262
rect 86 1258 90 1262
rect 102 1258 106 1262
rect 142 1258 146 1262
rect 6 1248 10 1252
rect 38 1248 42 1252
rect 22 1168 26 1172
rect 6 1148 10 1152
rect 78 1148 82 1152
rect 238 1298 242 1302
rect 286 1298 290 1302
rect 214 1278 218 1282
rect 238 1278 242 1282
rect 302 1288 306 1292
rect 206 1268 210 1272
rect 214 1268 218 1272
rect 342 1268 346 1272
rect 374 1268 378 1272
rect 262 1248 266 1252
rect 286 1248 290 1252
rect 302 1248 306 1252
rect 310 1248 314 1252
rect 174 1158 178 1162
rect 198 1158 202 1162
rect 262 1158 266 1162
rect 158 1148 162 1152
rect 286 1148 290 1152
rect 94 1138 98 1142
rect 54 1118 58 1122
rect 70 1118 74 1122
rect 14 1108 18 1112
rect 22 1098 26 1102
rect 174 1138 178 1142
rect 102 1118 106 1122
rect 166 1118 170 1122
rect 86 1108 90 1112
rect 86 1098 90 1102
rect 38 1088 42 1092
rect 70 1078 74 1082
rect 6 1068 10 1072
rect 22 1068 26 1072
rect 206 1138 210 1142
rect 230 1128 234 1132
rect 190 1108 194 1112
rect 206 1088 210 1092
rect 166 1068 170 1072
rect 102 1058 106 1062
rect 294 1098 298 1102
rect 318 1158 322 1162
rect 1002 1303 1006 1307
rect 1009 1303 1013 1307
rect 470 1278 474 1282
rect 478 1278 482 1282
rect 614 1278 618 1282
rect 1070 1278 1074 1282
rect 1094 1278 1098 1282
rect 1174 1278 1178 1282
rect 1214 1278 1218 1282
rect 1358 1278 1362 1282
rect 1478 1278 1482 1282
rect 430 1258 434 1262
rect 454 1258 458 1262
rect 462 1258 466 1262
rect 478 1258 482 1262
rect 414 1248 418 1252
rect 438 1238 442 1242
rect 462 1238 466 1242
rect 454 1228 458 1232
rect 398 1218 402 1222
rect 398 1148 402 1152
rect 398 1128 402 1132
rect 390 1118 394 1122
rect 406 1118 410 1122
rect 446 1148 450 1152
rect 430 1138 434 1142
rect 438 1128 442 1132
rect 430 1118 434 1122
rect 422 1098 426 1102
rect 358 1088 362 1092
rect 406 1088 410 1092
rect 438 1088 442 1092
rect 350 1078 354 1082
rect 526 1238 530 1242
rect 702 1268 706 1272
rect 806 1268 810 1272
rect 934 1268 938 1272
rect 982 1268 986 1272
rect 1062 1268 1066 1272
rect 582 1258 586 1262
rect 630 1248 634 1252
rect 598 1238 602 1242
rect 510 1228 514 1232
rect 534 1228 538 1232
rect 490 1203 494 1207
rect 497 1203 501 1207
rect 518 1158 522 1162
rect 526 1158 530 1162
rect 542 1158 546 1162
rect 550 1158 554 1162
rect 582 1158 586 1162
rect 654 1158 658 1162
rect 478 1148 482 1152
rect 598 1148 602 1152
rect 694 1208 698 1212
rect 678 1148 682 1152
rect 470 1138 474 1142
rect 502 1138 506 1142
rect 550 1138 554 1142
rect 566 1138 570 1142
rect 558 1128 562 1132
rect 606 1128 610 1132
rect 614 1128 618 1132
rect 502 1088 506 1092
rect 366 1068 370 1072
rect 430 1068 434 1072
rect 486 1068 490 1072
rect 550 1068 554 1072
rect 230 1058 234 1062
rect 22 1048 26 1052
rect 46 1048 50 1052
rect 214 1048 218 1052
rect 38 968 42 972
rect 6 948 10 952
rect 22 948 26 952
rect 94 958 98 962
rect 134 958 138 962
rect 198 958 202 962
rect 54 948 58 952
rect 86 940 90 944
rect 30 928 34 932
rect 6 868 10 872
rect 22 868 26 872
rect 46 868 50 872
rect 22 848 26 852
rect 30 848 34 852
rect 110 888 114 892
rect 102 878 106 882
rect 118 878 122 882
rect 134 878 138 882
rect 158 878 162 882
rect 182 878 186 882
rect 78 858 82 862
rect 118 858 122 862
rect 78 848 82 852
rect 102 848 106 852
rect 86 838 90 842
rect 190 858 194 862
rect 174 848 178 852
rect 30 828 34 832
rect 70 828 74 832
rect 158 828 162 832
rect 6 778 10 782
rect 38 748 42 752
rect 46 748 50 752
rect 118 748 122 752
rect 54 738 58 742
rect 150 758 154 762
rect 174 758 178 762
rect 182 758 186 762
rect 134 748 138 752
rect 22 728 26 732
rect 94 728 98 732
rect 110 728 114 732
rect 126 728 130 732
rect 22 718 26 722
rect 38 718 42 722
rect 30 688 34 692
rect 46 688 50 692
rect 446 1058 450 1062
rect 462 1058 466 1062
rect 534 1058 538 1062
rect 366 1048 370 1052
rect 446 1048 450 1052
rect 262 948 266 952
rect 318 968 322 972
rect 302 938 306 942
rect 214 888 218 892
rect 214 858 218 862
rect 278 848 282 852
rect 270 838 274 842
rect 310 838 314 842
rect 230 747 234 751
rect 166 738 170 742
rect 206 728 210 732
rect 214 708 218 712
rect 174 698 178 702
rect 286 768 290 772
rect 542 1038 546 1042
rect 490 1003 494 1007
rect 497 1003 501 1007
rect 358 998 362 1002
rect 374 998 378 1002
rect 582 1048 586 1052
rect 566 1038 570 1042
rect 438 958 442 962
rect 390 948 394 952
rect 406 948 410 952
rect 462 948 466 952
rect 374 928 378 932
rect 382 928 386 932
rect 406 928 410 932
rect 366 918 370 922
rect 526 918 530 922
rect 502 908 506 912
rect 502 878 506 882
rect 406 868 410 872
rect 430 868 434 872
rect 486 858 490 862
rect 366 788 370 792
rect 342 748 346 752
rect 358 708 362 712
rect 126 688 130 692
rect 326 688 330 692
rect 46 678 50 682
rect 94 678 98 682
rect 22 668 26 672
rect 86 668 90 672
rect 102 668 106 672
rect 174 678 178 682
rect 286 678 290 682
rect 14 658 18 662
rect 150 658 154 662
rect 158 658 162 662
rect 238 658 242 662
rect 150 648 154 652
rect 230 648 234 652
rect 318 658 322 662
rect 190 638 194 642
rect 294 638 298 642
rect 38 558 42 562
rect 110 588 114 592
rect 126 588 130 592
rect 318 588 322 592
rect 86 558 90 562
rect 30 528 34 532
rect 86 528 90 532
rect 6 478 10 482
rect 46 478 50 482
rect 246 568 250 572
rect 294 558 298 562
rect 350 558 354 562
rect 238 548 242 552
rect 262 548 266 552
rect 326 538 330 542
rect 150 528 154 532
rect 174 528 178 532
rect 118 518 122 522
rect 182 518 186 522
rect 166 478 170 482
rect 6 468 10 472
rect 110 468 114 472
rect 62 458 66 462
rect 94 458 98 462
rect 142 458 146 462
rect 22 448 26 452
rect 30 448 34 452
rect 78 448 82 452
rect 198 448 202 452
rect 182 418 186 422
rect 70 368 74 372
rect 6 358 10 362
rect 62 358 66 362
rect 94 358 98 362
rect 158 358 162 362
rect 30 348 34 352
rect 214 528 218 532
rect 246 528 250 532
rect 262 528 266 532
rect 334 528 338 532
rect 414 758 418 762
rect 518 848 522 852
rect 490 803 494 807
rect 497 803 501 807
rect 430 748 434 752
rect 374 738 378 742
rect 526 738 530 742
rect 398 688 402 692
rect 486 718 490 722
rect 494 678 498 682
rect 430 668 434 672
rect 398 548 402 552
rect 510 648 514 652
rect 478 628 482 632
rect 422 538 426 542
rect 382 528 386 532
rect 526 608 530 612
rect 490 603 494 607
rect 497 603 501 607
rect 662 1058 666 1062
rect 614 1048 618 1052
rect 662 1038 666 1042
rect 654 1018 658 1022
rect 582 958 586 962
rect 606 958 610 962
rect 566 938 570 942
rect 550 928 554 932
rect 590 928 594 932
rect 670 1018 674 1022
rect 606 938 610 942
rect 638 938 642 942
rect 638 928 642 932
rect 646 928 650 932
rect 630 918 634 922
rect 574 878 578 882
rect 582 878 586 882
rect 550 618 554 622
rect 638 868 642 872
rect 590 818 594 822
rect 638 818 642 822
rect 574 788 578 792
rect 574 778 578 782
rect 662 898 666 902
rect 686 1048 690 1052
rect 790 1258 794 1262
rect 862 1258 866 1262
rect 758 1238 762 1242
rect 726 1228 730 1232
rect 790 1218 794 1222
rect 886 1258 890 1262
rect 902 1258 906 1262
rect 926 1258 930 1262
rect 918 1238 922 1242
rect 878 1198 882 1202
rect 958 1228 962 1232
rect 966 1228 970 1232
rect 942 1218 946 1222
rect 926 1198 930 1202
rect 862 1168 866 1172
rect 894 1168 898 1172
rect 910 1168 914 1172
rect 814 1158 818 1162
rect 878 1158 882 1162
rect 726 1118 730 1122
rect 782 1108 786 1112
rect 854 1138 858 1142
rect 822 1118 826 1122
rect 814 1068 818 1072
rect 774 1058 778 1062
rect 798 1058 802 1062
rect 750 1038 754 1042
rect 702 1018 706 1022
rect 742 978 746 982
rect 750 958 754 962
rect 686 948 690 952
rect 710 948 714 952
rect 702 938 706 942
rect 734 948 738 952
rect 726 938 730 942
rect 678 928 682 932
rect 718 928 722 932
rect 718 908 722 912
rect 750 938 754 942
rect 758 928 762 932
rect 902 1158 906 1162
rect 902 1138 906 1142
rect 894 1108 898 1112
rect 958 1208 962 1212
rect 974 1208 978 1212
rect 982 1198 986 1202
rect 1014 1258 1018 1262
rect 1046 1258 1050 1262
rect 934 1188 938 1192
rect 942 1188 946 1192
rect 1006 1188 1010 1192
rect 950 1178 954 1182
rect 958 1158 962 1162
rect 990 1158 994 1162
rect 966 1138 970 1142
rect 982 1138 986 1142
rect 998 1128 1002 1132
rect 934 1118 938 1122
rect 1062 1238 1066 1242
rect 1046 1178 1050 1182
rect 1070 1188 1074 1192
rect 1094 1258 1098 1262
rect 1118 1258 1122 1262
rect 1126 1258 1130 1262
rect 1110 1208 1114 1212
rect 1126 1188 1130 1192
rect 1190 1178 1194 1182
rect 1182 1168 1186 1172
rect 1222 1258 1226 1262
rect 1262 1248 1266 1252
rect 1374 1268 1378 1272
rect 1318 1258 1322 1262
rect 1350 1258 1354 1262
rect 1254 1238 1258 1242
rect 1286 1238 1290 1242
rect 1310 1238 1314 1242
rect 1238 1228 1242 1232
rect 1326 1218 1330 1222
rect 1350 1228 1354 1232
rect 1390 1248 1394 1252
rect 1382 1238 1386 1242
rect 1374 1218 1378 1222
rect 1334 1208 1338 1212
rect 1366 1208 1370 1212
rect 1350 1198 1354 1202
rect 1254 1188 1258 1192
rect 1222 1178 1226 1182
rect 1246 1178 1250 1182
rect 1278 1178 1282 1182
rect 1214 1168 1218 1172
rect 1262 1168 1266 1172
rect 1126 1138 1130 1142
rect 1238 1138 1242 1142
rect 1014 1118 1018 1122
rect 1070 1118 1074 1122
rect 974 1108 978 1112
rect 1002 1103 1006 1107
rect 1009 1103 1013 1107
rect 926 1088 930 1092
rect 1014 1088 1018 1092
rect 878 1078 882 1082
rect 918 1078 922 1082
rect 838 1058 842 1062
rect 822 1018 826 1022
rect 830 1008 834 1012
rect 870 1058 874 1062
rect 910 1058 914 1062
rect 894 1048 898 1052
rect 854 1038 858 1042
rect 886 1038 890 1042
rect 886 1028 890 1032
rect 870 998 874 1002
rect 902 1028 906 1032
rect 950 1058 954 1062
rect 958 1048 962 1052
rect 966 1048 970 1052
rect 942 1028 946 1032
rect 990 1068 994 1072
rect 982 1058 986 1062
rect 974 1038 978 1042
rect 966 1018 970 1022
rect 854 988 858 992
rect 1358 1178 1362 1182
rect 1398 1218 1402 1222
rect 1398 1208 1402 1212
rect 1390 1158 1394 1162
rect 1350 1148 1354 1152
rect 1374 1148 1378 1152
rect 1382 1148 1386 1152
rect 1414 1198 1418 1202
rect 1454 1188 1458 1192
rect 1422 1168 1426 1172
rect 1438 1168 1442 1172
rect 1414 1158 1418 1162
rect 1198 1128 1202 1132
rect 1254 1128 1258 1132
rect 1286 1128 1290 1132
rect 1182 1118 1186 1122
rect 1150 1078 1154 1082
rect 1126 1068 1130 1072
rect 1070 1058 1074 1062
rect 1182 1058 1186 1062
rect 1198 1058 1202 1062
rect 1046 1048 1050 1052
rect 1078 1048 1082 1052
rect 1118 1048 1122 1052
rect 1150 1048 1154 1052
rect 838 978 842 982
rect 958 978 962 982
rect 998 978 1002 982
rect 798 968 802 972
rect 854 968 858 972
rect 870 968 874 972
rect 934 968 938 972
rect 942 968 946 972
rect 822 958 826 962
rect 838 948 842 952
rect 686 898 690 902
rect 678 888 682 892
rect 758 888 762 892
rect 654 878 658 882
rect 654 868 658 872
rect 678 868 682 872
rect 718 858 722 862
rect 710 848 714 852
rect 582 768 586 772
rect 606 768 610 772
rect 622 768 626 772
rect 638 768 642 772
rect 622 758 626 762
rect 646 748 650 752
rect 686 838 690 842
rect 686 768 690 772
rect 678 758 682 762
rect 702 758 706 762
rect 670 748 674 752
rect 638 738 642 742
rect 662 738 666 742
rect 630 728 634 732
rect 590 718 594 722
rect 598 718 602 722
rect 646 728 650 732
rect 590 708 594 712
rect 582 598 586 602
rect 558 588 562 592
rect 478 578 482 582
rect 542 578 546 582
rect 438 518 442 522
rect 462 518 466 522
rect 430 488 434 492
rect 606 688 610 692
rect 622 658 626 662
rect 606 648 610 652
rect 614 648 618 652
rect 502 568 506 572
rect 558 568 562 572
rect 590 568 594 572
rect 662 678 666 682
rect 646 668 650 672
rect 678 668 682 672
rect 686 668 690 672
rect 654 658 658 662
rect 694 658 698 662
rect 646 648 650 652
rect 742 858 746 862
rect 734 838 738 842
rect 726 768 730 772
rect 718 758 722 762
rect 710 748 714 752
rect 774 858 778 862
rect 766 838 770 842
rect 790 768 794 772
rect 830 938 834 942
rect 846 918 850 922
rect 806 868 810 872
rect 830 868 834 872
rect 822 848 826 852
rect 862 908 866 912
rect 862 898 866 902
rect 1014 968 1018 972
rect 894 958 898 962
rect 966 958 970 962
rect 982 958 986 962
rect 878 948 882 952
rect 934 948 938 952
rect 902 918 906 922
rect 918 918 922 922
rect 902 908 906 912
rect 918 888 922 892
rect 862 878 866 882
rect 846 778 850 782
rect 854 768 858 772
rect 798 758 802 762
rect 838 758 842 762
rect 750 748 754 752
rect 766 748 770 752
rect 798 748 802 752
rect 702 628 706 632
rect 638 618 642 622
rect 670 618 674 622
rect 702 598 706 602
rect 614 568 618 572
rect 630 568 634 572
rect 662 568 666 572
rect 526 558 530 562
rect 542 558 546 562
rect 590 558 594 562
rect 510 548 514 552
rect 542 548 546 552
rect 606 548 610 552
rect 534 538 538 542
rect 566 538 570 542
rect 582 538 586 542
rect 622 538 626 542
rect 638 548 642 552
rect 686 548 690 552
rect 734 708 738 712
rect 734 678 738 682
rect 718 638 722 642
rect 726 608 730 612
rect 910 868 914 872
rect 894 858 898 862
rect 894 838 898 842
rect 886 818 890 822
rect 870 808 874 812
rect 854 748 858 752
rect 918 768 922 772
rect 990 938 994 942
rect 1014 938 1018 942
rect 942 928 946 932
rect 974 908 978 912
rect 966 888 970 892
rect 966 878 970 882
rect 1002 903 1006 907
rect 1009 903 1013 907
rect 942 868 946 872
rect 982 868 986 872
rect 1014 868 1018 872
rect 958 858 962 862
rect 974 858 978 862
rect 942 828 946 832
rect 966 818 970 822
rect 950 808 954 812
rect 966 798 970 802
rect 958 758 962 762
rect 918 748 922 752
rect 934 748 938 752
rect 790 738 794 742
rect 862 738 866 742
rect 870 738 874 742
rect 894 738 898 742
rect 742 568 746 572
rect 742 558 746 562
rect 630 528 634 532
rect 654 538 658 542
rect 750 538 754 542
rect 822 708 826 712
rect 774 678 778 682
rect 846 698 850 702
rect 838 678 842 682
rect 790 668 794 672
rect 766 658 770 662
rect 798 658 802 662
rect 774 648 778 652
rect 806 648 810 652
rect 790 638 794 642
rect 806 638 810 642
rect 798 628 802 632
rect 774 618 778 622
rect 774 548 778 552
rect 854 678 858 682
rect 662 528 666 532
rect 638 518 642 522
rect 582 508 586 512
rect 446 488 450 492
rect 630 498 634 502
rect 350 478 354 482
rect 398 478 402 482
rect 566 478 570 482
rect 606 478 610 482
rect 230 468 234 472
rect 422 468 426 472
rect 278 458 282 462
rect 318 458 322 462
rect 206 388 210 392
rect 222 388 226 392
rect 270 388 274 392
rect 214 358 218 362
rect 110 348 114 352
rect 126 348 130 352
rect 182 348 186 352
rect 54 338 58 342
rect 94 338 98 342
rect 310 338 314 342
rect 350 458 354 462
rect 382 458 386 462
rect 390 458 394 462
rect 382 448 386 452
rect 406 448 410 452
rect 430 448 434 452
rect 334 438 338 442
rect 374 358 378 362
rect 422 358 426 362
rect 478 468 482 472
rect 454 458 458 462
rect 470 458 474 462
rect 486 458 490 462
rect 462 448 466 452
rect 622 458 626 462
rect 694 498 698 502
rect 662 468 666 472
rect 678 458 682 462
rect 694 458 698 462
rect 702 448 706 452
rect 702 438 706 442
rect 526 428 530 432
rect 598 428 602 432
rect 646 428 650 432
rect 490 403 494 407
rect 497 403 501 407
rect 638 408 642 412
rect 454 368 458 372
rect 486 358 490 362
rect 670 358 674 362
rect 470 338 474 342
rect 398 288 402 292
rect 406 288 410 292
rect 334 278 338 282
rect 14 268 18 272
rect 38 268 42 272
rect 70 268 74 272
rect 206 268 210 272
rect 214 268 218 272
rect 310 268 314 272
rect 94 248 98 252
rect 158 248 162 252
rect 238 258 242 262
rect 62 238 66 242
rect 142 238 146 242
rect 86 228 90 232
rect 54 148 58 152
rect 94 218 98 222
rect 166 148 170 152
rect 198 138 202 142
rect 110 128 114 132
rect 134 128 138 132
rect 118 118 122 122
rect 142 118 146 122
rect 150 118 154 122
rect 102 78 106 82
rect 70 68 74 72
rect 302 258 306 262
rect 262 238 266 242
rect 350 248 354 252
rect 446 218 450 222
rect 422 168 426 172
rect 542 328 546 332
rect 518 288 522 292
rect 510 278 514 282
rect 478 268 482 272
rect 490 203 494 207
rect 497 203 501 207
rect 470 158 474 162
rect 494 158 498 162
rect 414 148 418 152
rect 446 148 450 152
rect 486 148 490 152
rect 254 118 258 122
rect 438 138 442 142
rect 454 128 458 132
rect 462 128 466 132
rect 606 338 610 342
rect 654 328 658 332
rect 630 288 634 292
rect 582 278 586 282
rect 710 308 714 312
rect 574 258 578 262
rect 558 238 562 242
rect 614 168 618 172
rect 606 148 610 152
rect 542 138 546 142
rect 574 138 578 142
rect 246 88 250 92
rect 270 88 274 92
rect 694 188 698 192
rect 702 178 706 182
rect 638 138 642 142
rect 646 138 650 142
rect 166 78 170 82
rect 302 78 306 82
rect 334 78 338 82
rect 350 78 354 82
rect 446 78 450 82
rect 542 78 546 82
rect 118 68 122 72
rect 270 68 274 72
rect 78 58 82 62
rect 166 58 170 62
rect 198 58 202 62
rect 6 48 10 52
rect 70 48 74 52
rect 86 38 90 42
rect 182 48 186 52
rect 270 58 274 62
rect 550 68 554 72
rect 318 58 322 62
rect 326 58 330 62
rect 342 58 346 62
rect 278 48 282 52
rect 398 58 402 62
rect 438 59 442 63
rect 798 528 802 532
rect 814 528 818 532
rect 726 518 730 522
rect 782 518 786 522
rect 838 518 842 522
rect 734 478 738 482
rect 822 508 826 512
rect 806 488 810 492
rect 814 478 818 482
rect 750 458 754 462
rect 734 448 738 452
rect 750 438 754 442
rect 774 458 778 462
rect 830 498 834 502
rect 846 478 850 482
rect 790 448 794 452
rect 806 448 810 452
rect 822 448 826 452
rect 798 418 802 422
rect 814 378 818 382
rect 750 358 754 362
rect 766 358 770 362
rect 806 358 810 362
rect 726 338 730 342
rect 734 338 738 342
rect 718 288 722 292
rect 742 318 746 322
rect 726 158 730 162
rect 734 148 738 152
rect 806 348 810 352
rect 766 338 770 342
rect 774 328 778 332
rect 750 138 754 142
rect 718 78 722 82
rect 790 318 794 322
rect 774 278 778 282
rect 766 178 770 182
rect 766 168 770 172
rect 870 548 874 552
rect 902 728 906 732
rect 910 728 914 732
rect 910 698 914 702
rect 934 688 938 692
rect 910 678 914 682
rect 894 668 898 672
rect 918 668 922 672
rect 942 668 946 672
rect 902 648 906 652
rect 934 648 938 652
rect 886 628 890 632
rect 910 588 914 592
rect 926 588 930 592
rect 902 568 906 572
rect 870 538 874 542
rect 878 538 882 542
rect 1030 1038 1034 1042
rect 1046 1038 1050 1042
rect 1038 1018 1042 1022
rect 1062 1038 1066 1042
rect 1086 1038 1090 1042
rect 1110 1038 1114 1042
rect 1054 1008 1058 1012
rect 1110 1028 1114 1032
rect 1030 978 1034 982
rect 1086 978 1090 982
rect 1126 978 1130 982
rect 1094 968 1098 972
rect 1118 968 1122 972
rect 1054 958 1058 962
rect 1118 958 1122 962
rect 1030 938 1034 942
rect 1038 928 1042 932
rect 1038 918 1042 922
rect 1038 908 1042 912
rect 1022 858 1026 862
rect 990 788 994 792
rect 998 778 1002 782
rect 1014 838 1018 842
rect 1006 768 1010 772
rect 982 758 986 762
rect 1022 768 1026 772
rect 990 738 994 742
rect 982 728 986 732
rect 1070 948 1074 952
rect 1062 938 1066 942
rect 1102 938 1106 942
rect 1190 1048 1194 1052
rect 1174 1038 1178 1042
rect 1214 1038 1218 1042
rect 1438 1138 1442 1142
rect 1302 1118 1306 1122
rect 1342 1118 1346 1122
rect 1414 1118 1418 1122
rect 1446 1118 1450 1122
rect 1366 1088 1370 1092
rect 1406 1088 1410 1092
rect 1422 1088 1426 1092
rect 1334 1078 1338 1082
rect 1286 1068 1290 1072
rect 1278 1058 1282 1062
rect 1294 1058 1298 1062
rect 1254 1048 1258 1052
rect 1270 1038 1274 1042
rect 1166 1028 1170 1032
rect 1198 1028 1202 1032
rect 1230 1028 1234 1032
rect 1246 1028 1250 1032
rect 1174 1018 1178 1022
rect 1166 958 1170 962
rect 1190 968 1194 972
rect 1118 948 1122 952
rect 1150 948 1154 952
rect 1070 928 1074 932
rect 1046 888 1050 892
rect 1110 888 1114 892
rect 1070 878 1074 882
rect 1102 878 1106 882
rect 1062 858 1066 862
rect 1054 838 1058 842
rect 1094 858 1098 862
rect 1110 858 1114 862
rect 1246 1008 1250 1012
rect 1238 978 1242 982
rect 1214 958 1218 962
rect 1214 948 1218 952
rect 1166 938 1170 942
rect 1190 938 1194 942
rect 1278 998 1282 1002
rect 1270 978 1274 982
rect 1254 968 1258 972
rect 1286 968 1290 972
rect 1246 948 1250 952
rect 1270 948 1274 952
rect 1198 928 1202 932
rect 1206 928 1210 932
rect 1230 928 1234 932
rect 1142 908 1146 912
rect 1126 868 1130 872
rect 1166 878 1170 882
rect 1174 878 1178 882
rect 1150 868 1154 872
rect 1086 848 1090 852
rect 1110 848 1114 852
rect 1078 768 1082 772
rect 1302 1008 1306 1012
rect 1414 1078 1418 1082
rect 1430 1068 1434 1072
rect 1326 1058 1330 1062
rect 1342 1028 1346 1032
rect 1318 988 1322 992
rect 1310 978 1314 982
rect 1310 968 1314 972
rect 1326 968 1330 972
rect 1462 1158 1466 1162
rect 1486 1158 1490 1162
rect 1462 1118 1466 1122
rect 1470 1118 1474 1122
rect 1454 1078 1458 1082
rect 1446 1058 1450 1062
rect 1350 998 1354 1002
rect 1366 1048 1370 1052
rect 1382 1048 1386 1052
rect 1422 1048 1426 1052
rect 1358 988 1362 992
rect 1310 958 1314 962
rect 1374 998 1378 1002
rect 1406 998 1410 1002
rect 1390 988 1394 992
rect 1310 948 1314 952
rect 1334 948 1338 952
rect 1366 948 1370 952
rect 1390 948 1394 952
rect 1342 938 1346 942
rect 1286 918 1290 922
rect 1294 918 1298 922
rect 1318 918 1322 922
rect 1238 888 1242 892
rect 1214 878 1218 882
rect 1182 848 1186 852
rect 1182 838 1186 842
rect 1134 828 1138 832
rect 1174 828 1178 832
rect 1118 798 1122 802
rect 1206 828 1210 832
rect 1262 868 1266 872
rect 1270 858 1274 862
rect 1302 858 1306 862
rect 1318 868 1322 872
rect 1350 858 1354 862
rect 1238 848 1242 852
rect 1310 848 1314 852
rect 1486 1098 1490 1102
rect 1494 1098 1498 1102
rect 1494 1078 1498 1082
rect 1478 1068 1482 1072
rect 1502 1068 1506 1072
rect 1462 1058 1466 1062
rect 1486 1048 1490 1052
rect 1438 968 1442 972
rect 1478 968 1482 972
rect 1510 1048 1514 1052
rect 1486 948 1490 952
rect 1502 948 1506 952
rect 1462 938 1466 942
rect 1470 938 1474 942
rect 1430 928 1434 932
rect 1438 898 1442 902
rect 1430 888 1434 892
rect 1414 878 1418 882
rect 1438 878 1442 882
rect 1446 878 1450 882
rect 1406 868 1410 872
rect 1382 858 1386 862
rect 1430 858 1434 862
rect 1478 888 1482 892
rect 1462 868 1466 872
rect 1486 878 1490 882
rect 1454 858 1458 862
rect 1390 848 1394 852
rect 1438 848 1442 852
rect 1462 848 1466 852
rect 1302 838 1306 842
rect 1334 838 1338 842
rect 1366 838 1370 842
rect 1398 838 1402 842
rect 1462 838 1466 842
rect 1470 838 1474 842
rect 1246 828 1250 832
rect 1302 828 1306 832
rect 1350 828 1354 832
rect 1214 818 1218 822
rect 1118 768 1122 772
rect 1142 778 1146 782
rect 1190 778 1194 782
rect 1206 778 1210 782
rect 1262 778 1266 782
rect 1358 808 1362 812
rect 1414 808 1418 812
rect 1390 798 1394 802
rect 1390 788 1394 792
rect 1398 778 1402 782
rect 1150 768 1154 772
rect 1134 758 1138 762
rect 1166 758 1170 762
rect 1078 748 1082 752
rect 1110 748 1114 752
rect 1126 748 1130 752
rect 1070 738 1074 742
rect 1086 738 1090 742
rect 1222 768 1226 772
rect 1238 768 1242 772
rect 1278 768 1282 772
rect 1286 768 1290 772
rect 1390 768 1394 772
rect 1422 768 1426 772
rect 1222 748 1226 752
rect 1270 758 1274 762
rect 1310 758 1314 762
rect 1382 758 1386 762
rect 1206 738 1210 742
rect 1246 738 1250 742
rect 1286 738 1290 742
rect 1046 728 1050 732
rect 1062 728 1066 732
rect 1110 728 1114 732
rect 1126 728 1130 732
rect 1198 728 1202 732
rect 1206 728 1210 732
rect 1246 728 1250 732
rect 1262 728 1266 732
rect 1014 718 1018 722
rect 1002 703 1006 707
rect 1009 703 1013 707
rect 990 688 994 692
rect 1030 688 1034 692
rect 1078 678 1082 682
rect 1126 678 1130 682
rect 1150 678 1154 682
rect 1062 668 1066 672
rect 1198 688 1202 692
rect 1190 678 1194 682
rect 1262 688 1266 692
rect 1214 678 1218 682
rect 1246 678 1250 682
rect 1206 668 1210 672
rect 1214 668 1218 672
rect 1222 668 1226 672
rect 1254 668 1258 672
rect 1038 658 1042 662
rect 1102 658 1106 662
rect 1158 658 1162 662
rect 1030 648 1034 652
rect 1158 648 1162 652
rect 1174 648 1178 652
rect 1190 648 1194 652
rect 1230 658 1234 662
rect 1286 658 1290 662
rect 1406 758 1410 762
rect 1382 748 1386 752
rect 1310 658 1314 662
rect 1286 648 1290 652
rect 1294 648 1298 652
rect 1318 648 1322 652
rect 1142 638 1146 642
rect 966 618 970 622
rect 982 608 986 612
rect 942 568 946 572
rect 1086 608 1090 612
rect 1062 588 1066 592
rect 1094 588 1098 592
rect 1126 588 1130 592
rect 1038 578 1042 582
rect 1078 578 1082 582
rect 990 568 994 572
rect 1062 568 1066 572
rect 1046 558 1050 562
rect 1070 558 1074 562
rect 942 548 946 552
rect 958 548 962 552
rect 990 548 994 552
rect 1014 548 1018 552
rect 974 538 978 542
rect 1014 538 1018 542
rect 1022 538 1026 542
rect 878 528 882 532
rect 918 528 922 532
rect 966 528 970 532
rect 870 518 874 522
rect 902 518 906 522
rect 870 508 874 512
rect 926 508 930 512
rect 966 508 970 512
rect 870 478 874 482
rect 942 478 946 482
rect 1014 528 1018 532
rect 1038 528 1042 532
rect 982 498 986 502
rect 982 488 986 492
rect 1002 503 1006 507
rect 1009 503 1013 507
rect 1102 578 1106 582
rect 1118 568 1122 572
rect 1134 578 1138 582
rect 1150 578 1154 582
rect 1150 568 1154 572
rect 1166 568 1170 572
rect 1142 548 1146 552
rect 1078 528 1082 532
rect 1054 518 1058 522
rect 1110 508 1114 512
rect 1118 498 1122 502
rect 1030 488 1034 492
rect 1078 488 1082 492
rect 990 478 994 482
rect 1110 478 1114 482
rect 862 468 866 472
rect 902 468 906 472
rect 974 468 978 472
rect 1006 468 1010 472
rect 1070 468 1074 472
rect 1374 728 1378 732
rect 1446 768 1450 772
rect 1462 768 1466 772
rect 1486 828 1490 832
rect 1478 768 1482 772
rect 1502 938 1506 942
rect 1510 898 1514 902
rect 1478 758 1482 762
rect 1494 758 1498 762
rect 1454 748 1458 752
rect 1486 748 1490 752
rect 1502 738 1506 742
rect 1430 688 1434 692
rect 1382 678 1386 682
rect 1334 658 1338 662
rect 1350 648 1354 652
rect 1422 658 1426 662
rect 1438 658 1442 662
rect 1374 648 1378 652
rect 1430 648 1434 652
rect 1334 638 1338 642
rect 1366 638 1370 642
rect 1334 628 1338 632
rect 1406 628 1410 632
rect 1326 598 1330 602
rect 1310 588 1314 592
rect 1238 578 1242 582
rect 1302 578 1306 582
rect 1182 568 1186 572
rect 1246 568 1250 572
rect 1278 568 1282 572
rect 1310 568 1314 572
rect 1230 558 1234 562
rect 1254 558 1258 562
rect 1174 548 1178 552
rect 1230 548 1234 552
rect 1174 538 1178 542
rect 1190 538 1194 542
rect 1270 548 1274 552
rect 1286 548 1290 552
rect 1294 538 1298 542
rect 1198 528 1202 532
rect 1222 528 1226 532
rect 1230 528 1234 532
rect 1278 528 1282 532
rect 1286 528 1290 532
rect 1198 518 1202 522
rect 1150 488 1154 492
rect 1150 478 1154 482
rect 878 458 882 462
rect 894 458 898 462
rect 1102 458 1106 462
rect 854 448 858 452
rect 838 428 842 432
rect 838 378 842 382
rect 886 358 890 362
rect 854 348 858 352
rect 862 348 866 352
rect 910 448 914 452
rect 934 448 938 452
rect 958 448 962 452
rect 910 358 914 362
rect 926 348 930 352
rect 878 338 882 342
rect 894 338 898 342
rect 918 338 922 342
rect 934 338 938 342
rect 830 328 834 332
rect 870 328 874 332
rect 862 298 866 302
rect 830 268 834 272
rect 854 268 858 272
rect 870 268 874 272
rect 910 328 914 332
rect 894 318 898 322
rect 934 318 938 322
rect 902 288 906 292
rect 958 308 962 312
rect 942 278 946 282
rect 950 268 954 272
rect 838 258 842 262
rect 1038 448 1042 452
rect 1054 448 1058 452
rect 974 358 978 362
rect 974 328 978 332
rect 1054 348 1058 352
rect 1094 348 1098 352
rect 1150 468 1154 472
rect 1166 468 1170 472
rect 1262 518 1266 522
rect 1270 508 1274 512
rect 1238 488 1242 492
rect 1206 468 1210 472
rect 1174 458 1178 462
rect 1190 458 1194 462
rect 1134 368 1138 372
rect 1126 358 1130 362
rect 1182 358 1186 362
rect 1118 348 1122 352
rect 1150 348 1154 352
rect 1030 338 1034 342
rect 1070 338 1074 342
rect 1110 338 1114 342
rect 1002 303 1006 307
rect 1009 303 1013 307
rect 1030 288 1034 292
rect 1070 318 1074 322
rect 1102 308 1106 312
rect 1110 288 1114 292
rect 974 258 978 262
rect 910 248 914 252
rect 822 188 826 192
rect 1006 278 1010 282
rect 1046 278 1050 282
rect 990 258 994 262
rect 1126 328 1130 332
rect 1254 468 1258 472
rect 1222 438 1226 442
rect 1262 438 1266 442
rect 1246 358 1250 362
rect 1358 578 1362 582
rect 1350 568 1354 572
rect 1374 568 1378 572
rect 1342 548 1346 552
rect 1326 518 1330 522
rect 1334 508 1338 512
rect 1318 488 1322 492
rect 1310 468 1314 472
rect 1382 528 1386 532
rect 1350 488 1354 492
rect 1374 488 1378 492
rect 1382 468 1386 472
rect 1366 458 1370 462
rect 1374 458 1378 462
rect 1326 438 1330 442
rect 1358 438 1362 442
rect 1358 418 1362 422
rect 1310 358 1314 362
rect 1230 348 1234 352
rect 1262 348 1266 352
rect 1278 348 1282 352
rect 1134 308 1138 312
rect 1142 298 1146 302
rect 1126 278 1130 282
rect 1030 268 1034 272
rect 1078 268 1082 272
rect 1118 268 1122 272
rect 1150 288 1154 292
rect 1166 288 1170 292
rect 1062 258 1066 262
rect 1094 258 1098 262
rect 1102 258 1106 262
rect 998 248 1002 252
rect 1046 248 1050 252
rect 1070 248 1074 252
rect 1054 198 1058 202
rect 1046 178 1050 182
rect 926 168 930 172
rect 950 168 954 172
rect 1022 168 1026 172
rect 1030 168 1034 172
rect 854 158 858 162
rect 774 148 778 152
rect 838 148 842 152
rect 766 138 770 142
rect 822 138 826 142
rect 1094 178 1098 182
rect 934 158 938 162
rect 950 158 954 162
rect 1062 158 1066 162
rect 1070 158 1074 162
rect 1094 158 1098 162
rect 942 148 946 152
rect 1054 148 1058 152
rect 798 128 802 132
rect 830 128 834 132
rect 854 128 858 132
rect 902 138 906 142
rect 918 138 922 142
rect 974 138 978 142
rect 1022 138 1026 142
rect 1110 188 1114 192
rect 1102 148 1106 152
rect 1118 168 1122 172
rect 1190 278 1194 282
rect 1214 278 1218 282
rect 1174 268 1178 272
rect 1198 268 1202 272
rect 1238 338 1242 342
rect 1254 338 1258 342
rect 1254 328 1258 332
rect 1190 238 1194 242
rect 1158 198 1162 202
rect 1254 278 1258 282
rect 1270 278 1274 282
rect 1254 268 1258 272
rect 1246 188 1250 192
rect 1222 168 1226 172
rect 1262 168 1266 172
rect 1150 158 1154 162
rect 1158 148 1162 152
rect 1254 158 1258 162
rect 1238 148 1242 152
rect 1334 358 1338 362
rect 1294 288 1298 292
rect 1310 288 1314 292
rect 1366 358 1370 362
rect 1342 328 1346 332
rect 1334 278 1338 282
rect 1286 268 1290 272
rect 1318 268 1322 272
rect 1366 268 1370 272
rect 1294 258 1298 262
rect 1310 258 1314 262
rect 1334 258 1338 262
rect 1318 248 1322 252
rect 1286 218 1290 222
rect 1270 148 1274 152
rect 1326 148 1330 152
rect 1382 418 1386 422
rect 1398 598 1402 602
rect 1430 588 1434 592
rect 1462 678 1466 682
rect 1454 648 1458 652
rect 1470 588 1474 592
rect 1446 578 1450 582
rect 1486 578 1490 582
rect 1510 598 1514 602
rect 1478 548 1482 552
rect 1494 548 1498 552
rect 1398 538 1402 542
rect 1406 538 1410 542
rect 1486 538 1490 542
rect 1398 468 1402 472
rect 1454 488 1458 492
rect 1454 468 1458 472
rect 1486 468 1490 472
rect 1414 458 1418 462
rect 1470 458 1474 462
rect 1398 448 1402 452
rect 1430 448 1434 452
rect 1446 438 1450 442
rect 1470 438 1474 442
rect 1390 358 1394 362
rect 1462 368 1466 372
rect 1382 348 1386 352
rect 1430 348 1434 352
rect 1438 348 1442 352
rect 1390 338 1394 342
rect 1406 338 1410 342
rect 1422 328 1426 332
rect 1414 318 1418 322
rect 1446 308 1450 312
rect 1438 268 1442 272
rect 1470 308 1474 312
rect 1470 298 1474 302
rect 1454 268 1458 272
rect 1382 258 1386 262
rect 1374 248 1378 252
rect 1350 238 1354 242
rect 1366 228 1370 232
rect 1398 248 1402 252
rect 1430 248 1434 252
rect 1462 248 1466 252
rect 1414 238 1418 242
rect 1446 238 1450 242
rect 1406 228 1410 232
rect 1390 218 1394 222
rect 1374 158 1378 162
rect 1078 138 1082 142
rect 1142 138 1146 142
rect 1206 138 1210 142
rect 1262 138 1266 142
rect 966 128 970 132
rect 1230 128 1234 132
rect 878 118 882 122
rect 1214 118 1218 122
rect 758 68 762 72
rect 798 68 802 72
rect 490 3 494 7
rect 497 3 501 7
rect 878 68 882 72
rect 910 68 914 72
rect 862 58 866 62
rect 1002 103 1006 107
rect 1009 103 1013 107
rect 998 78 1002 82
rect 1118 78 1122 82
rect 1014 68 1018 72
rect 1238 78 1242 82
rect 1358 78 1362 82
rect 982 58 986 62
rect 1486 268 1490 272
rect 1478 178 1482 182
rect 1486 158 1490 162
rect 1462 148 1466 152
rect 1478 138 1482 142
rect 1454 128 1458 132
rect 1470 128 1474 132
rect 1502 138 1506 142
rect 1390 58 1394 62
rect 1422 58 1426 62
rect 1470 58 1474 62
<< metal3 >>
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1014 1303 1016 1307
rect 242 1298 286 1301
rect 178 1288 302 1291
rect 18 1278 54 1281
rect 218 1278 238 1281
rect 474 1278 478 1281
rect 1074 1278 1094 1281
rect -26 1271 -22 1272
rect -26 1268 22 1271
rect 114 1268 166 1271
rect 210 1268 214 1271
rect 614 1271 617 1278
rect 378 1268 617 1271
rect 706 1268 806 1271
rect 810 1268 870 1271
rect 986 1268 1062 1271
rect 1174 1271 1177 1278
rect 1066 1268 1177 1271
rect 1214 1271 1217 1278
rect 1214 1268 1350 1271
rect 1358 1271 1361 1278
rect 1478 1272 1481 1278
rect 1358 1268 1374 1271
rect 66 1258 70 1261
rect 90 1258 102 1261
rect 342 1261 345 1268
rect 146 1258 345 1261
rect 434 1258 449 1261
rect 458 1258 462 1261
rect 586 1258 633 1261
rect -26 1251 -22 1252
rect -26 1248 6 1251
rect 10 1248 38 1251
rect 266 1248 286 1251
rect 290 1248 302 1251
rect 314 1248 350 1251
rect 354 1248 414 1251
rect 446 1251 449 1258
rect 478 1251 481 1258
rect 418 1248 441 1251
rect 446 1248 481 1251
rect 630 1252 633 1258
rect 866 1258 886 1261
rect 906 1258 926 1261
rect 934 1261 937 1268
rect 934 1258 1014 1261
rect 1050 1258 1094 1261
rect 1130 1258 1134 1261
rect 1226 1258 1318 1261
rect 1322 1258 1350 1261
rect 790 1251 793 1258
rect 1118 1251 1121 1258
rect 790 1248 1121 1251
rect 1266 1248 1270 1251
rect 1354 1248 1390 1251
rect 438 1242 441 1248
rect 466 1238 526 1241
rect 530 1238 598 1241
rect 762 1238 918 1241
rect 922 1238 1062 1241
rect 1258 1238 1286 1241
rect 1314 1238 1382 1241
rect 458 1228 510 1231
rect 514 1228 534 1231
rect 730 1228 958 1231
rect 1242 1228 1350 1231
rect 402 1218 406 1221
rect 694 1218 742 1221
rect 794 1218 942 1221
rect 966 1221 969 1228
rect 966 1218 1326 1221
rect 1330 1218 1374 1221
rect 1402 1218 1470 1221
rect 694 1212 697 1218
rect 962 1208 974 1211
rect 1114 1208 1334 1211
rect 1338 1208 1366 1211
rect 1370 1208 1398 1211
rect 488 1203 490 1207
rect 494 1203 497 1207
rect 502 1203 504 1207
rect 882 1198 926 1201
rect 930 1198 982 1201
rect 1354 1198 1414 1201
rect 946 1188 1006 1191
rect 1010 1188 1070 1191
rect 1258 1188 1454 1191
rect 934 1181 937 1188
rect 934 1178 950 1181
rect 954 1178 1046 1181
rect 1126 1181 1129 1188
rect 1126 1178 1190 1181
rect 1194 1178 1222 1181
rect 1226 1178 1246 1181
rect 1250 1178 1278 1181
rect -26 1171 -22 1172
rect -26 1168 22 1171
rect 866 1168 894 1171
rect 914 1168 1182 1171
rect 1186 1168 1214 1171
rect 1218 1168 1262 1171
rect 1358 1171 1361 1178
rect 1358 1168 1422 1171
rect 1442 1168 1454 1171
rect 178 1158 198 1161
rect 266 1158 318 1161
rect 522 1158 526 1161
rect 546 1158 550 1161
rect 554 1158 582 1161
rect 818 1158 878 1161
rect 906 1158 958 1161
rect 962 1158 990 1161
rect 1394 1158 1414 1161
rect 1418 1158 1462 1161
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 10 1148 78 1151
rect 402 1148 414 1151
rect 450 1148 478 1151
rect 654 1151 657 1158
rect 1486 1152 1489 1158
rect 602 1148 657 1151
rect 682 1148 1262 1151
rect 1266 1148 1350 1151
rect 1378 1148 1382 1151
rect 158 1141 161 1148
rect 98 1138 174 1141
rect 286 1141 289 1148
rect 210 1138 289 1141
rect 434 1138 470 1141
rect 474 1138 502 1141
rect 554 1138 566 1141
rect 858 1138 862 1141
rect 906 1138 966 1141
rect 986 1138 1126 1141
rect 1242 1138 1438 1141
rect 62 1128 230 1131
rect 402 1128 438 1131
rect 562 1128 606 1131
rect 610 1128 614 1131
rect 966 1131 969 1138
rect 1198 1132 1201 1138
rect 966 1128 998 1131
rect 1258 1128 1286 1131
rect 1466 1128 1473 1131
rect 62 1121 65 1128
rect 1470 1122 1473 1128
rect 58 1118 65 1121
rect 74 1118 102 1121
rect 106 1118 166 1121
rect 394 1118 406 1121
rect 418 1118 430 1121
rect 730 1118 822 1121
rect 938 1118 1014 1121
rect 1018 1118 1070 1121
rect 1186 1118 1302 1121
rect 1346 1118 1414 1121
rect 1450 1118 1462 1121
rect 18 1108 86 1111
rect 90 1108 190 1111
rect 786 1108 894 1111
rect 898 1108 974 1111
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1014 1103 1016 1107
rect 26 1098 86 1101
rect 298 1098 414 1101
rect 426 1098 438 1101
rect 1402 1098 1486 1101
rect 1494 1092 1497 1098
rect 210 1088 358 1091
rect 410 1088 438 1091
rect 442 1088 502 1091
rect 930 1088 1014 1091
rect 1202 1088 1366 1091
rect 1410 1088 1422 1091
rect 38 1081 41 1088
rect 38 1078 70 1081
rect 882 1078 918 1081
rect 978 1078 1150 1081
rect 1338 1078 1414 1081
rect 1458 1078 1494 1081
rect 350 1072 353 1078
rect -26 1071 -22 1072
rect -26 1068 6 1071
rect 10 1068 22 1071
rect 370 1068 430 1071
rect 490 1068 550 1071
rect 818 1068 982 1071
rect 994 1068 1126 1071
rect 1290 1068 1430 1071
rect 1482 1068 1502 1071
rect 166 1061 169 1068
rect 982 1062 985 1068
rect 166 1058 230 1061
rect 450 1058 462 1061
rect 538 1058 585 1061
rect -26 1051 -22 1052
rect -26 1048 22 1051
rect 26 1048 46 1051
rect 102 1051 105 1058
rect 582 1052 585 1058
rect 618 1058 662 1061
rect 778 1058 798 1061
rect 842 1058 870 1061
rect 914 1058 950 1061
rect 1074 1058 1182 1061
rect 1186 1058 1198 1061
rect 1202 1058 1278 1061
rect 1298 1058 1326 1061
rect 1382 1058 1446 1061
rect 1466 1058 1470 1061
rect 614 1052 617 1058
rect 686 1052 689 1058
rect 1382 1052 1385 1058
rect 102 1048 214 1051
rect 370 1048 446 1051
rect 898 1048 902 1051
rect 906 1048 958 1051
rect 970 1048 1046 1051
rect 1050 1048 1070 1051
rect 1082 1048 1118 1051
rect 1194 1048 1254 1051
rect 1258 1048 1366 1051
rect 1426 1048 1462 1051
rect 1490 1048 1510 1051
rect 546 1038 566 1041
rect 666 1038 750 1041
rect 858 1038 886 1041
rect 978 1038 1030 1041
rect 1050 1038 1062 1041
rect 1090 1038 1110 1041
rect 1150 1041 1153 1048
rect 1150 1038 1174 1041
rect 1178 1038 1214 1041
rect 1218 1038 1270 1041
rect 878 1028 886 1031
rect 890 1028 902 1031
rect 906 1028 942 1031
rect 1102 1028 1110 1031
rect 1114 1028 1166 1031
rect 1202 1028 1230 1031
rect 1242 1028 1246 1031
rect 1250 1028 1342 1031
rect 650 1018 654 1021
rect 674 1018 702 1021
rect 826 1018 966 1021
rect 1042 1018 1174 1021
rect 834 1008 1054 1011
rect 1250 1008 1302 1011
rect 488 1003 490 1007
rect 494 1003 497 1007
rect 502 1003 504 1007
rect 1054 1002 1057 1008
rect 362 998 374 1001
rect 874 998 1046 1001
rect 1282 998 1350 1001
rect 1354 998 1374 1001
rect 1378 998 1406 1001
rect 846 988 854 991
rect 858 988 1318 991
rect 1322 988 1358 991
rect 1362 988 1390 991
rect 746 978 838 981
rect 842 978 958 981
rect 1002 978 1030 981
rect 1034 978 1086 981
rect 1130 978 1238 981
rect 1242 978 1270 981
rect 1274 978 1310 981
rect -26 971 -22 972
rect -26 968 38 971
rect 42 968 318 971
rect 790 968 798 971
rect 802 968 854 971
rect 874 968 934 971
rect 938 968 942 971
rect 946 968 1014 971
rect 1098 968 1118 971
rect 1122 968 1190 971
rect 1290 968 1310 971
rect 1314 968 1326 971
rect 1442 968 1470 971
rect 1474 968 1478 971
rect 98 958 110 961
rect 586 958 606 961
rect 754 958 822 961
rect 890 958 894 961
rect 970 958 982 961
rect 986 958 1054 961
rect 1058 958 1118 961
rect 1170 958 1214 961
rect 1254 961 1257 968
rect 1254 958 1310 961
rect -26 951 -22 952
rect -26 948 6 951
rect 26 948 54 951
rect 134 951 137 958
rect 198 951 201 958
rect 438 952 441 958
rect 1502 952 1505 958
rect 134 948 201 951
rect 266 948 390 951
rect 394 948 406 951
rect 466 948 614 951
rect 690 948 710 951
rect 714 948 734 951
rect 842 948 878 951
rect 938 948 1070 951
rect 1122 948 1150 951
rect 1218 948 1246 951
rect 1250 948 1270 951
rect 1314 948 1334 951
rect 1370 948 1390 951
rect 1458 948 1486 951
rect 30 940 86 941
rect 30 938 89 940
rect 298 938 302 941
rect 570 938 606 941
rect 642 938 702 941
rect 706 938 726 941
rect 754 938 830 941
rect 986 938 990 941
rect 1018 938 1030 941
rect 1066 938 1070 941
rect 1074 938 1102 941
rect 1170 938 1190 941
rect 1346 938 1433 941
rect 1466 938 1470 941
rect 1482 938 1502 941
rect 30 932 33 938
rect 942 932 945 938
rect 1430 932 1433 938
rect 378 928 382 931
rect 410 928 550 931
rect 554 928 590 931
rect 642 928 646 931
rect 682 928 718 931
rect 722 928 758 931
rect 1042 928 1070 931
rect 1074 928 1198 931
rect 1210 928 1230 931
rect 370 918 526 921
rect 634 918 686 921
rect 850 918 902 921
rect 922 918 1038 921
rect 1290 918 1294 921
rect 1298 918 1318 921
rect 482 908 502 911
rect 722 908 862 911
rect 906 908 974 911
rect 1042 908 1142 911
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1014 903 1016 907
rect 666 898 686 901
rect 858 898 862 901
rect 1442 898 1478 901
rect 1510 892 1513 898
rect 114 888 214 891
rect 654 888 678 891
rect 762 888 918 891
rect 970 888 1046 891
rect 1114 888 1238 891
rect 1434 888 1454 891
rect 1458 888 1478 891
rect 654 882 657 888
rect 106 878 118 881
rect 122 878 134 881
rect 150 878 158 881
rect 162 878 182 881
rect 578 878 582 881
rect 866 878 966 881
rect 1074 878 1102 881
rect 1178 878 1214 881
rect 1418 878 1438 881
rect 1450 878 1486 881
rect -26 871 -22 872
rect -26 868 6 871
rect 18 868 22 871
rect 26 868 46 871
rect 50 868 406 871
rect 502 871 505 878
rect 434 868 505 871
rect 642 868 654 871
rect 682 868 806 871
rect 826 868 830 871
rect 834 868 910 871
rect 946 868 958 871
rect 986 868 1014 871
rect 1018 868 1070 871
rect 1074 868 1126 871
rect 1130 868 1150 871
rect 1166 871 1169 878
rect 1166 868 1262 871
rect 1322 868 1326 871
rect 1382 868 1406 871
rect 1450 868 1462 871
rect 718 862 721 868
rect 1382 862 1385 868
rect 82 858 118 861
rect 194 858 214 861
rect 490 858 521 861
rect 746 858 774 861
rect 898 858 958 861
rect 962 858 974 861
rect 978 858 1022 861
rect 1026 858 1062 861
rect 1066 858 1094 861
rect 1114 858 1270 861
rect 1306 858 1350 861
rect 1354 858 1382 861
rect 1394 858 1430 861
rect 1434 858 1454 861
rect 518 852 521 858
rect 1390 852 1393 858
rect -26 851 -22 852
rect -26 848 14 851
rect 26 848 30 851
rect 82 848 102 851
rect 178 848 278 851
rect 714 848 822 851
rect 906 848 1086 851
rect 1114 848 1182 851
rect 1242 848 1310 851
rect 1442 848 1462 851
rect 30 838 86 841
rect 274 838 310 841
rect 650 838 686 841
rect 690 838 734 841
rect 746 838 766 841
rect 770 838 894 841
rect 1018 838 1054 841
rect 1186 838 1302 841
rect 1306 838 1334 841
rect 1370 838 1398 841
rect 1458 838 1462 841
rect 1474 838 1494 841
rect 30 832 33 838
rect 74 828 158 831
rect 886 828 918 831
rect 922 828 942 831
rect 946 828 1134 831
rect 1138 828 1174 831
rect 1210 828 1246 831
rect 1306 828 1350 831
rect 1354 828 1486 831
rect 886 822 889 828
rect 586 818 590 821
rect 594 818 638 821
rect 958 818 966 821
rect 970 818 1214 821
rect 874 808 942 811
rect 946 808 950 811
rect 1362 808 1414 811
rect 488 803 490 807
rect 494 803 497 807
rect 502 803 504 807
rect 890 798 966 801
rect 970 798 1118 801
rect 1394 798 1398 801
rect 370 788 574 791
rect 898 788 990 791
rect -26 781 -22 782
rect -26 778 6 781
rect 578 778 846 781
rect 1002 778 1142 781
rect 1146 778 1190 781
rect 1194 778 1206 781
rect 1250 778 1262 781
rect 1390 781 1393 788
rect 1354 778 1393 781
rect 1402 778 1457 781
rect 1454 772 1457 778
rect 586 768 590 771
rect 610 768 622 771
rect 642 768 646 771
rect 690 768 726 771
rect 730 768 790 771
rect 794 768 854 771
rect 922 768 1006 771
rect 1010 768 1022 771
rect 1082 768 1118 771
rect 1122 768 1150 771
rect 1226 768 1238 771
rect 1242 768 1278 771
rect 1394 768 1398 771
rect 1426 768 1446 771
rect 1458 768 1462 771
rect 1466 768 1478 771
rect -26 761 -22 762
rect -26 758 121 761
rect 154 758 174 761
rect 178 758 182 761
rect 286 761 289 768
rect 286 758 414 761
rect 626 758 678 761
rect 682 758 702 761
rect 722 758 798 761
rect 842 758 958 761
rect 962 758 982 761
rect 1138 758 1166 761
rect 1286 761 1289 768
rect 1286 758 1310 761
rect 1386 758 1406 761
rect 1410 758 1438 761
rect 1482 758 1494 761
rect 118 752 121 758
rect 42 748 46 751
rect 122 748 134 751
rect 138 748 230 751
rect 346 748 430 751
rect 594 748 646 751
rect 650 748 670 751
rect 674 748 710 751
rect 742 748 750 751
rect 754 748 766 751
rect 770 748 798 751
rect 858 748 918 751
rect 1082 748 1110 751
rect 1130 748 1222 751
rect 1270 751 1273 758
rect 1226 748 1273 751
rect 1386 748 1390 751
rect 1402 748 1454 751
rect 934 742 937 748
rect 1206 742 1209 748
rect -26 741 -22 742
rect -26 738 54 741
rect 378 738 526 741
rect 642 738 662 741
rect 794 738 862 741
rect 874 738 894 741
rect 994 738 1070 741
rect 1074 738 1086 741
rect 1250 738 1286 741
rect 1486 741 1489 748
rect 1474 738 1489 741
rect 10 728 22 731
rect 98 728 110 731
rect 166 731 169 738
rect 130 728 169 731
rect 206 732 209 738
rect 902 732 905 738
rect 1374 732 1377 738
rect 1502 732 1505 738
rect 634 728 646 731
rect 914 728 982 731
rect 1050 728 1062 731
rect 1066 728 1110 731
rect 1130 728 1198 731
rect 1210 728 1246 731
rect 1250 728 1262 731
rect 14 718 22 721
rect 26 718 38 721
rect 490 718 590 721
rect 602 718 878 721
rect 942 718 1014 721
rect 218 708 302 711
rect 362 708 406 711
rect 594 708 734 711
rect 942 711 945 718
rect 826 708 945 711
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1014 703 1016 707
rect -26 701 -22 702
rect -26 698 14 701
rect 850 698 910 701
rect 174 692 177 698
rect -26 688 30 691
rect 50 688 126 691
rect 330 688 398 691
rect 586 688 606 691
rect 994 688 1030 691
rect 1202 688 1262 691
rect 1434 688 1462 691
rect -26 682 -23 688
rect -26 678 -22 682
rect 18 678 46 681
rect 98 678 174 681
rect 666 678 734 681
rect 770 678 774 681
rect 842 678 854 681
rect 858 678 910 681
rect 934 681 937 688
rect 934 678 1073 681
rect 1082 678 1126 681
rect 1154 678 1190 681
rect 1194 678 1214 681
rect 1254 678 1382 681
rect 26 668 86 671
rect 106 668 110 671
rect 286 671 289 678
rect 114 668 289 671
rect 494 671 497 678
rect 918 672 921 678
rect 434 668 497 671
rect 642 668 646 671
rect 650 668 678 671
rect 690 668 790 671
rect 890 668 894 671
rect 946 668 1062 671
rect 1070 671 1073 678
rect 1246 672 1249 678
rect 1254 672 1257 678
rect 1070 668 1206 671
rect 1226 668 1246 671
rect 1462 671 1465 678
rect 1378 668 1465 671
rect -26 661 -22 662
rect -26 658 6 661
rect 10 658 14 661
rect 86 661 89 668
rect 86 658 150 661
rect 162 658 238 661
rect 322 658 513 661
rect 626 658 654 661
rect 658 658 694 661
rect 698 658 766 661
rect 802 658 998 661
rect 1042 658 1102 661
rect 1214 661 1217 668
rect 1162 658 1230 661
rect 1234 658 1286 661
rect 1314 658 1334 661
rect 1426 658 1438 661
rect 510 652 513 658
rect 154 648 158 651
rect 162 648 230 651
rect 610 648 614 651
rect 650 648 766 651
rect 778 648 806 651
rect 906 648 934 651
rect 938 648 1030 651
rect 1162 648 1174 651
rect 1178 648 1185 651
rect 1194 648 1198 651
rect 1250 648 1286 651
rect 1298 648 1302 651
rect 1322 648 1350 651
rect 1354 648 1374 651
rect 1434 648 1454 651
rect 194 638 294 641
rect 722 638 790 641
rect 810 638 1142 641
rect 1146 638 1334 641
rect 1338 638 1366 641
rect 482 628 702 631
rect 706 628 798 631
rect 802 628 886 631
rect 1338 628 1406 631
rect 554 618 638 621
rect 642 618 670 621
rect 778 618 966 621
rect 530 608 726 611
rect 986 608 1086 611
rect 488 603 490 607
rect 494 603 497 607
rect 502 603 504 607
rect 514 598 582 601
rect 706 598 1326 601
rect 1330 598 1398 601
rect 1402 598 1510 601
rect 114 588 126 591
rect 310 588 318 591
rect 322 588 558 591
rect 914 588 926 591
rect 930 588 1062 591
rect 1098 588 1126 591
rect 1130 588 1310 591
rect 1434 588 1470 591
rect 482 578 542 581
rect 1082 578 1102 581
rect 1106 578 1134 581
rect 1138 578 1150 581
rect 1242 578 1289 581
rect 1294 578 1302 581
rect 1306 578 1358 581
rect 1362 578 1446 581
rect 506 568 558 571
rect 562 568 590 571
rect 594 568 614 571
rect 658 568 662 571
rect 666 568 742 571
rect 906 568 942 571
rect 946 568 990 571
rect 1038 571 1041 578
rect 1038 568 1062 571
rect 1122 568 1150 571
rect 1154 568 1166 571
rect 1186 568 1246 571
rect 1250 568 1278 571
rect 1286 571 1289 578
rect 1286 568 1310 571
rect 1486 571 1489 578
rect 1378 568 1489 571
rect 246 561 249 568
rect 246 558 294 561
rect 298 558 350 561
rect 530 558 542 561
rect 630 561 633 568
rect 1350 562 1353 568
rect 594 558 742 561
rect 942 558 1046 561
rect 1074 558 1230 561
rect 1234 558 1254 561
rect 38 551 41 558
rect 86 551 89 558
rect 942 552 945 558
rect 1478 552 1481 558
rect 38 548 89 551
rect 242 548 262 551
rect 266 548 278 551
rect 514 548 542 551
rect 610 548 638 551
rect 690 548 774 551
rect 874 548 886 551
rect 962 548 990 551
rect 1018 548 1142 551
rect 1178 548 1230 551
rect 1234 548 1270 551
rect 1290 548 1342 551
rect 1482 548 1494 551
rect 398 541 401 548
rect 330 538 401 541
rect 426 538 534 541
rect 570 538 582 541
rect 586 538 590 541
rect 626 538 654 541
rect 754 538 870 541
rect 882 538 974 541
rect 986 538 1014 541
rect 1026 538 1030 541
rect 1178 538 1190 541
rect 1230 538 1294 541
rect 1402 538 1406 541
rect 1466 538 1486 541
rect 1230 532 1233 538
rect 34 528 86 531
rect 154 528 174 531
rect 218 528 246 531
rect 250 528 262 531
rect 338 528 382 531
rect 634 528 662 531
rect 802 528 806 531
rect 810 528 814 531
rect 870 528 878 531
rect 882 528 918 531
rect 970 528 1014 531
rect 1018 528 1038 531
rect 1082 528 1198 531
rect 1226 528 1230 531
rect 1262 528 1278 531
rect 1282 528 1286 531
rect 1378 528 1382 531
rect 870 522 873 528
rect 1262 522 1265 528
rect 122 518 182 521
rect 186 518 206 521
rect 442 518 462 521
rect 642 518 726 521
rect 786 518 838 521
rect 842 518 854 521
rect 894 518 902 521
rect 906 518 958 521
rect 966 518 1046 521
rect 1058 518 1198 521
rect 1314 518 1326 521
rect 966 512 969 518
rect 586 508 822 511
rect 874 508 918 511
rect 930 508 934 511
rect 1114 508 1270 511
rect 1274 508 1334 511
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1014 503 1016 507
rect 634 498 694 501
rect 834 498 982 501
rect 1034 498 1118 501
rect 594 488 806 491
rect 814 488 974 491
rect 986 488 1030 491
rect 1034 488 1078 491
rect 1154 488 1238 491
rect 1242 488 1318 491
rect 1322 488 1350 491
rect 1458 488 1470 491
rect 10 478 46 481
rect 354 478 382 481
rect 430 481 433 488
rect 402 478 433 481
rect 446 482 449 488
rect 814 482 817 488
rect 1374 482 1377 488
rect 610 478 734 481
rect 866 478 870 481
rect 890 478 942 481
rect 946 478 982 481
rect 994 478 1110 481
rect 1114 478 1150 481
rect -26 471 -22 472
rect -26 468 6 471
rect 166 471 169 478
rect 114 468 169 471
rect 426 468 478 471
rect 566 471 569 478
rect 482 468 569 471
rect 846 471 849 478
rect 666 468 849 471
rect 866 468 902 471
rect 978 468 1006 471
rect 1010 468 1070 471
rect 1170 468 1174 471
rect 1178 468 1206 471
rect 1258 468 1310 471
rect 1386 468 1398 471
rect 1402 468 1454 471
rect 1458 468 1486 471
rect 66 458 94 461
rect 230 461 233 468
rect 146 458 201 461
rect 230 458 278 461
rect 322 458 350 461
rect 354 458 382 461
rect 394 458 454 461
rect 474 458 486 461
rect 618 458 622 461
rect 626 458 678 461
rect 698 458 750 461
rect 778 458 878 461
rect 898 458 966 461
rect 986 458 1102 461
rect 1150 461 1153 468
rect 1150 458 1174 461
rect 1178 458 1190 461
rect 1370 458 1374 461
rect 1378 458 1414 461
rect 1418 458 1470 461
rect 198 452 201 458
rect -26 451 -22 452
rect -26 448 22 451
rect 34 448 78 451
rect 386 448 406 451
rect 434 448 462 451
rect 706 448 734 451
rect 782 448 790 451
rect 794 448 806 451
rect 826 448 854 451
rect 858 448 910 451
rect 914 448 934 451
rect 962 448 1038 451
rect 1042 448 1054 451
rect 1402 448 1430 451
rect 1446 442 1449 448
rect 10 438 334 441
rect 338 438 702 441
rect 754 438 1222 441
rect 1226 438 1262 441
rect 1266 438 1326 441
rect 1330 438 1358 441
rect 1450 438 1470 441
rect 530 428 598 431
rect 650 428 838 431
rect 842 428 878 431
rect 178 418 182 421
rect 802 418 862 421
rect 1362 418 1374 421
rect 1378 418 1382 421
rect 642 408 654 411
rect 488 403 490 407
rect 494 403 497 407
rect 502 403 504 407
rect 210 388 222 391
rect 274 388 278 391
rect 810 378 814 381
rect 818 378 838 381
rect 882 368 1134 371
rect -26 361 -22 362
rect -26 358 6 361
rect 10 358 62 361
rect 70 361 73 368
rect 70 358 94 361
rect 162 358 214 361
rect 454 361 457 368
rect 1462 362 1465 368
rect 426 358 486 361
rect 754 358 766 361
rect 770 358 806 361
rect 858 358 886 361
rect 914 358 974 361
rect 1130 358 1182 361
rect 1250 358 1310 361
rect 1370 358 1390 361
rect 34 348 110 351
rect 130 348 182 351
rect 374 351 377 358
rect 670 351 673 358
rect 374 348 673 351
rect 810 348 854 351
rect 858 348 862 351
rect 930 348 937 351
rect 1058 348 1094 351
rect 1122 348 1150 351
rect 1234 348 1262 351
rect 1266 348 1278 351
rect 1334 351 1337 358
rect 1334 348 1382 351
rect 1434 348 1438 351
rect 934 342 937 348
rect -26 341 -22 342
rect -26 338 54 341
rect 58 338 94 341
rect 98 338 310 341
rect 474 338 545 341
rect 610 338 657 341
rect 730 338 734 341
rect 770 338 878 341
rect 898 338 918 341
rect 1034 338 1070 341
rect 1074 338 1110 341
rect 1242 338 1254 341
rect 1394 338 1406 341
rect 542 332 545 338
rect 654 332 657 338
rect 778 328 822 331
rect 834 328 870 331
rect 874 328 897 331
rect 914 328 974 331
rect 1070 328 1126 331
rect 1346 328 1422 331
rect 894 322 897 328
rect 1070 322 1073 328
rect 1254 322 1257 328
rect 746 318 790 321
rect 938 318 1070 321
rect 1258 318 1414 321
rect 714 308 902 311
rect 906 308 958 311
rect 1106 308 1134 311
rect 1450 308 1470 311
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1014 303 1016 307
rect 850 298 862 301
rect 1110 298 1142 301
rect 1474 298 1510 301
rect 1110 292 1113 298
rect 402 288 406 291
rect 514 288 518 291
rect 634 288 718 291
rect 722 288 894 291
rect 898 288 902 291
rect 1034 288 1110 291
rect 1154 288 1166 291
rect 1298 288 1310 291
rect 514 278 582 281
rect 854 278 942 281
rect 946 278 1006 281
rect 1010 278 1046 281
rect 1130 278 1190 281
rect 1218 278 1254 281
rect 1274 278 1334 281
rect -26 271 -22 272
rect -26 268 6 271
rect 10 268 14 271
rect 42 268 70 271
rect 210 268 214 271
rect 218 268 310 271
rect 334 271 337 278
rect 314 268 337 271
rect 774 271 777 278
rect 854 272 857 278
rect 774 268 830 271
rect 954 268 1030 271
rect 1082 268 1118 271
rect 1178 268 1198 271
rect 1202 268 1254 271
rect 1258 268 1286 271
rect 1314 268 1318 271
rect 1322 268 1366 271
rect 1442 268 1454 271
rect 238 262 241 268
rect 94 258 161 261
rect 478 261 481 268
rect 306 258 353 261
rect 478 258 574 261
rect 870 261 873 268
rect 842 258 873 261
rect 978 258 990 261
rect 1066 258 1094 261
rect 1106 258 1294 261
rect 1314 258 1334 261
rect 1338 258 1382 261
rect 1486 261 1489 268
rect 1442 258 1489 261
rect 94 252 97 258
rect 158 252 161 258
rect 350 252 353 258
rect 882 248 910 251
rect 1002 248 1046 251
rect 1050 248 1070 251
rect 1322 248 1374 251
rect 1402 248 1430 251
rect 1458 248 1462 251
rect 66 238 142 241
rect 266 238 558 241
rect 1194 238 1350 241
rect 1418 238 1446 241
rect 90 228 158 231
rect 1370 228 1406 231
rect 98 218 446 221
rect 1290 218 1390 221
rect 488 203 490 207
rect 494 203 497 207
rect 502 203 504 207
rect 1058 198 1158 201
rect 698 188 822 191
rect 1046 188 1110 191
rect 1114 188 1246 191
rect 1466 188 1481 191
rect 1046 182 1049 188
rect 1478 182 1481 188
rect 706 178 766 181
rect 618 168 729 171
rect 422 161 425 168
rect 726 162 729 168
rect 930 168 950 171
rect 1026 168 1030 171
rect 1094 171 1097 178
rect 1094 168 1118 171
rect 1226 168 1262 171
rect 422 158 470 161
rect 474 158 494 161
rect 766 161 769 168
rect 1486 162 1489 168
rect 766 158 854 161
rect 938 158 950 161
rect 954 158 1062 161
rect 1074 158 1094 161
rect 1098 158 1150 161
rect 1258 158 1262 161
rect -26 151 -22 152
rect -26 148 54 151
rect 170 148 201 151
rect 418 148 446 151
rect 490 148 545 151
rect 610 148 649 151
rect 738 148 774 151
rect 842 148 846 151
rect 902 148 942 151
rect 1058 148 1065 151
rect 1106 148 1158 151
rect 1242 148 1270 151
rect 1374 151 1377 158
rect 1330 148 1377 151
rect 1542 151 1546 152
rect 1466 148 1546 151
rect 198 142 201 148
rect 438 142 441 148
rect 542 142 545 148
rect 646 142 649 148
rect 902 142 905 148
rect 578 138 638 141
rect 754 138 766 141
rect 826 138 902 141
rect 978 138 1022 141
rect 1026 138 1078 141
rect 1082 138 1142 141
rect 1210 138 1262 141
rect 1482 138 1502 141
rect -26 131 -22 132
rect -26 128 110 131
rect 114 128 134 131
rect 458 128 462 131
rect 466 128 478 131
rect 834 128 854 131
rect 918 131 921 138
rect 918 128 966 131
rect 1214 128 1230 131
rect 1458 128 1470 131
rect 122 118 142 121
rect 154 118 254 121
rect 798 121 801 128
rect 1214 122 1217 128
rect 798 118 878 121
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1014 103 1016 107
rect 250 88 270 91
rect 106 78 166 81
rect 306 78 334 81
rect 338 78 350 81
rect 450 78 542 81
rect 1002 78 1118 81
rect 1122 78 1238 81
rect 1242 78 1358 81
rect 74 68 118 71
rect 274 68 550 71
rect 718 71 721 78
rect 718 68 758 71
rect 762 68 798 71
rect 998 71 1001 78
rect 914 68 1001 71
rect 82 58 166 61
rect 202 58 270 61
rect 322 58 326 61
rect 346 58 398 61
rect 402 59 438 61
rect 402 58 441 59
rect 878 61 881 68
rect 866 58 881 61
rect 1014 61 1017 68
rect 986 58 1017 61
rect 1394 58 1422 61
rect 1470 52 1473 58
rect -26 51 -22 52
rect -26 48 6 51
rect 74 48 89 51
rect 186 48 278 51
rect 86 42 89 48
rect 488 3 490 7
rect 494 3 497 7
rect 502 3 504 7
<< m4contact >>
rect 1002 1303 1006 1307
rect 1010 1303 1013 1307
rect 1013 1303 1014 1307
rect 870 1268 874 1272
rect 1350 1268 1354 1272
rect 1478 1268 1482 1272
rect 350 1248 354 1252
rect 1134 1258 1138 1262
rect 1270 1248 1274 1252
rect 1350 1248 1354 1252
rect 406 1218 410 1222
rect 742 1218 746 1222
rect 1470 1218 1474 1222
rect 490 1203 494 1207
rect 498 1203 501 1207
rect 501 1203 502 1207
rect 1454 1168 1458 1172
rect 414 1148 418 1152
rect 1262 1148 1266 1152
rect 1486 1148 1490 1152
rect 862 1138 866 1142
rect 1198 1138 1202 1142
rect 1462 1128 1466 1132
rect 414 1118 418 1122
rect 1002 1103 1006 1107
rect 1010 1103 1013 1107
rect 1013 1103 1014 1107
rect 414 1098 418 1102
rect 438 1098 442 1102
rect 1398 1098 1402 1102
rect 1198 1088 1202 1092
rect 1494 1088 1498 1092
rect 974 1078 978 1082
rect 350 1068 354 1072
rect 982 1068 986 1072
rect 614 1058 618 1062
rect 686 1058 690 1062
rect 1470 1058 1474 1062
rect 902 1048 906 1052
rect 1070 1048 1074 1052
rect 1462 1048 1466 1052
rect 1238 1028 1242 1032
rect 646 1018 650 1022
rect 490 1003 494 1007
rect 498 1003 501 1007
rect 501 1003 502 1007
rect 1046 998 1050 1002
rect 1054 998 1058 1002
rect 1470 968 1474 972
rect 110 958 114 962
rect 886 958 890 962
rect 1502 958 1506 962
rect 438 948 442 952
rect 614 948 618 952
rect 1454 948 1458 952
rect 294 938 298 942
rect 942 938 946 942
rect 982 938 986 942
rect 1070 938 1074 942
rect 1478 938 1482 942
rect 686 918 690 922
rect 478 908 482 912
rect 1002 903 1006 907
rect 1010 903 1013 907
rect 1013 903 1014 907
rect 854 898 858 902
rect 1478 898 1482 902
rect 1454 888 1458 892
rect 1510 888 1514 892
rect 14 868 18 872
rect 822 868 826 872
rect 958 868 962 872
rect 1070 868 1074 872
rect 1326 868 1330 872
rect 1446 868 1450 872
rect 1390 858 1394 862
rect 14 848 18 852
rect 902 848 906 852
rect 646 838 650 842
rect 742 838 746 842
rect 1054 838 1058 842
rect 1454 838 1458 842
rect 1494 838 1498 842
rect 918 828 922 832
rect 582 818 586 822
rect 942 808 946 812
rect 490 803 494 807
rect 498 803 501 807
rect 501 803 502 807
rect 886 798 890 802
rect 1398 798 1402 802
rect 894 788 898 792
rect 1246 778 1250 782
rect 1350 778 1354 782
rect 590 768 594 772
rect 646 768 650 772
rect 1398 768 1402 772
rect 1454 768 1458 772
rect 1438 758 1442 762
rect 590 748 594 752
rect 1390 748 1394 752
rect 1398 748 1402 752
rect 206 738 210 742
rect 902 738 906 742
rect 934 738 938 742
rect 1374 738 1378 742
rect 1470 738 1474 742
rect 6 728 10 732
rect 1502 728 1506 732
rect 878 718 882 722
rect 302 708 306 712
rect 406 708 410 712
rect 1002 703 1006 707
rect 1010 703 1013 707
rect 1013 703 1014 707
rect 14 698 18 702
rect 174 688 178 692
rect 582 688 586 692
rect 1462 688 1466 692
rect 14 678 18 682
rect 766 678 770 682
rect 918 678 922 682
rect 110 668 114 672
rect 638 668 642 672
rect 886 668 890 672
rect 1246 668 1250 672
rect 1374 668 1378 672
rect 6 658 10 662
rect 998 658 1002 662
rect 158 648 162 652
rect 766 648 770 652
rect 1198 648 1202 652
rect 1246 648 1250 652
rect 1302 648 1306 652
rect 490 603 494 607
rect 498 603 501 607
rect 501 603 502 607
rect 510 598 514 602
rect 654 568 658 572
rect 1350 558 1354 562
rect 1478 558 1482 562
rect 278 548 282 552
rect 886 548 890 552
rect 590 538 594 542
rect 982 538 986 542
rect 1030 538 1034 542
rect 1462 538 1466 542
rect 806 528 810 532
rect 1374 528 1378 532
rect 206 518 210 522
rect 854 518 858 522
rect 958 518 962 522
rect 1046 518 1050 522
rect 1310 518 1314 522
rect 918 508 922 512
rect 934 508 938 512
rect 1002 503 1006 507
rect 1010 503 1013 507
rect 1013 503 1014 507
rect 1030 498 1034 502
rect 590 488 594 492
rect 974 488 978 492
rect 1470 488 1474 492
rect 382 478 386 482
rect 446 478 450 482
rect 862 478 866 482
rect 886 478 890 482
rect 982 478 986 482
rect 1374 478 1378 482
rect 1174 468 1178 472
rect 614 458 618 462
rect 966 458 970 462
rect 982 458 986 462
rect 1446 448 1450 452
rect 6 438 10 442
rect 878 428 882 432
rect 174 418 178 422
rect 862 418 866 422
rect 1374 418 1378 422
rect 654 408 658 412
rect 490 403 494 407
rect 498 403 501 407
rect 501 403 502 407
rect 278 388 282 392
rect 806 378 810 382
rect 878 368 882 372
rect 854 358 858 362
rect 1462 358 1466 362
rect 822 328 826 332
rect 1254 318 1258 322
rect 902 308 906 312
rect 1002 303 1006 307
rect 1010 303 1013 307
rect 1013 303 1014 307
rect 846 298 850 302
rect 1510 298 1514 302
rect 510 288 514 292
rect 894 288 898 292
rect 6 268 10 272
rect 1310 268 1314 272
rect 1438 258 1442 262
rect 878 248 882 252
rect 1454 248 1458 252
rect 158 228 162 232
rect 490 203 494 207
rect 498 203 501 207
rect 501 203 502 207
rect 1462 188 1466 192
rect 1486 168 1490 172
rect 1262 158 1266 162
rect 846 148 850 152
rect 478 128 482 132
rect 1002 103 1006 107
rect 1010 103 1013 107
rect 1013 103 1014 107
rect 1470 48 1474 52
rect 490 3 494 7
rect 498 3 501 7
rect 501 3 502 7
<< metal4 >>
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1014 1303 1016 1307
rect 870 1262 873 1268
rect 1130 1258 1134 1261
rect 1350 1252 1353 1268
rect 1262 1248 1270 1251
rect 350 1072 353 1248
rect 14 852 17 868
rect 6 662 9 728
rect 14 682 17 698
rect 110 672 113 958
rect 298 938 305 941
rect 6 272 9 438
rect 158 232 161 648
rect 174 422 177 688
rect 206 522 209 738
rect 302 712 305 938
rect 406 712 409 1218
rect 488 1203 490 1207
rect 494 1203 497 1207
rect 502 1203 504 1207
rect 414 1122 417 1148
rect 414 1102 417 1118
rect 438 952 441 1098
rect 488 1003 490 1007
rect 494 1003 497 1007
rect 502 1003 504 1007
rect 614 952 617 1058
rect 278 392 281 548
rect 386 478 390 481
rect 442 478 446 481
rect 478 132 481 908
rect 488 803 490 807
rect 494 803 497 807
rect 502 803 504 807
rect 582 692 585 818
rect 590 752 593 768
rect 488 603 490 607
rect 494 603 497 607
rect 502 603 504 607
rect 488 403 490 407
rect 494 403 497 407
rect 502 403 504 407
rect 510 292 513 598
rect 590 542 593 748
rect 590 492 593 538
rect 614 462 617 948
rect 646 842 649 1018
rect 686 922 689 1058
rect 742 842 745 1218
rect 1262 1152 1265 1248
rect 854 1138 862 1141
rect 854 902 857 1138
rect 1198 1132 1201 1138
rect 638 768 646 771
rect 638 672 641 768
rect 766 652 769 678
rect 654 412 657 568
rect 806 382 809 528
rect 822 332 825 868
rect 878 722 881 1128
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1014 1103 1016 1107
rect 1198 1092 1201 1128
rect 886 802 889 958
rect 902 852 905 1048
rect 894 671 897 788
rect 890 668 897 671
rect 854 362 857 518
rect 886 482 889 548
rect 862 422 865 478
rect 878 372 881 428
rect 488 203 490 207
rect 494 203 497 207
rect 502 203 504 207
rect 846 152 849 298
rect 878 252 881 368
rect 894 292 897 668
rect 902 742 905 848
rect 902 312 905 738
rect 918 682 921 828
rect 942 812 945 938
rect 962 868 966 871
rect 974 861 977 1078
rect 982 942 985 1068
rect 1046 1002 1049 1028
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1014 903 1016 907
rect 966 858 977 861
rect 918 512 921 528
rect 934 512 937 738
rect 958 522 961 538
rect 966 462 969 858
rect 1054 842 1057 998
rect 1070 942 1073 1048
rect 1242 1028 1246 1031
rect 1070 872 1073 938
rect 1322 868 1326 871
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1014 703 1016 707
rect 1246 672 1249 778
rect 998 652 1001 658
rect 1246 652 1249 668
rect 1194 648 1198 651
rect 1298 648 1302 651
rect 1350 562 1353 778
rect 1390 752 1393 858
rect 1398 802 1401 1098
rect 1454 952 1457 1168
rect 1462 1052 1465 1128
rect 1470 1062 1473 1218
rect 1398 772 1401 798
rect 1398 752 1401 768
rect 1374 672 1377 738
rect 974 538 982 541
rect 1026 538 1030 541
rect 974 492 977 538
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1014 503 1016 507
rect 1030 502 1033 538
rect 1374 532 1377 668
rect 1378 528 1382 531
rect 982 462 985 478
rect 1046 472 1049 518
rect 1170 468 1174 471
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1014 303 1016 307
rect 1254 161 1257 318
rect 1310 272 1313 518
rect 1374 422 1377 478
rect 1438 262 1441 758
rect 1446 452 1449 868
rect 1454 842 1457 888
rect 1454 252 1457 768
rect 1470 742 1473 968
rect 1478 942 1481 1268
rect 1462 542 1465 688
rect 1478 562 1481 898
rect 1462 192 1465 358
rect 1254 158 1262 161
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1014 103 1016 107
rect 1470 52 1473 488
rect 1486 172 1489 1148
rect 1494 842 1497 1088
rect 1502 732 1505 958
rect 1510 302 1513 888
rect 488 3 490 7
rect 494 3 497 7
rect 502 3 504 7
<< m5contact >>
rect 1002 1303 1006 1307
rect 1009 1303 1010 1307
rect 1010 1303 1013 1307
rect 870 1258 874 1262
rect 1126 1258 1130 1262
rect 490 1203 494 1207
rect 497 1203 498 1207
rect 498 1203 501 1207
rect 490 1003 494 1007
rect 497 1003 498 1007
rect 498 1003 501 1007
rect 390 478 394 482
rect 438 478 442 482
rect 490 803 494 807
rect 497 803 498 807
rect 498 803 501 807
rect 490 603 494 607
rect 497 603 498 607
rect 498 603 501 607
rect 490 403 494 407
rect 497 403 498 407
rect 498 403 501 407
rect 878 1128 882 1132
rect 1198 1128 1202 1132
rect 1002 1103 1006 1107
rect 1009 1103 1010 1107
rect 1010 1103 1013 1107
rect 490 203 494 207
rect 497 203 498 207
rect 498 203 501 207
rect 966 868 970 872
rect 1046 1028 1050 1032
rect 1002 903 1006 907
rect 1009 903 1010 907
rect 1010 903 1013 907
rect 918 528 922 532
rect 958 538 962 542
rect 1246 1028 1250 1032
rect 1318 868 1322 872
rect 1002 703 1006 707
rect 1009 703 1010 707
rect 1010 703 1013 707
rect 998 648 1002 652
rect 1190 648 1194 652
rect 1294 648 1298 652
rect 1022 538 1026 542
rect 1002 503 1006 507
rect 1009 503 1010 507
rect 1010 503 1013 507
rect 1382 528 1386 532
rect 1046 468 1050 472
rect 1166 468 1170 472
rect 1002 303 1006 307
rect 1009 303 1010 307
rect 1010 303 1013 307
rect 1002 103 1006 107
rect 1009 103 1010 107
rect 1010 103 1013 107
rect 490 3 494 7
rect 497 3 498 7
rect 498 3 501 7
<< metal5 >>
rect 1006 1303 1009 1307
rect 1005 1302 1010 1303
rect 1015 1302 1016 1307
rect 874 1258 1126 1261
rect 494 1203 497 1207
rect 493 1202 498 1203
rect 503 1202 504 1207
rect 882 1128 1198 1131
rect 1006 1103 1009 1107
rect 1005 1102 1010 1103
rect 1015 1102 1016 1107
rect 1050 1028 1246 1031
rect 494 1003 497 1007
rect 493 1002 498 1003
rect 503 1002 504 1007
rect 1006 903 1009 907
rect 1005 902 1010 903
rect 1015 902 1016 907
rect 970 868 1318 871
rect 494 803 497 807
rect 493 802 498 803
rect 503 802 504 807
rect 1006 703 1009 707
rect 1005 702 1010 703
rect 1015 702 1016 707
rect 1002 648 1190 651
rect 1194 648 1294 651
rect 494 603 497 607
rect 493 602 498 603
rect 503 602 504 607
rect 962 538 1022 541
rect 922 528 1382 531
rect 1006 503 1009 507
rect 1005 502 1010 503
rect 1015 502 1016 507
rect 394 478 438 481
rect 1050 468 1166 471
rect 494 403 497 407
rect 493 402 498 403
rect 503 402 504 407
rect 1006 303 1009 307
rect 1005 302 1010 303
rect 1015 302 1016 307
rect 494 203 497 207
rect 493 202 498 203
rect 503 202 504 207
rect 1006 103 1009 107
rect 1005 102 1010 103
rect 1015 102 1016 107
rect 494 3 497 7
rect 493 2 498 3
rect 503 2 504 7
<< m6contact >>
rect 1000 1303 1002 1307
rect 1002 1303 1005 1307
rect 1010 1303 1013 1307
rect 1013 1303 1015 1307
rect 1000 1302 1005 1303
rect 1010 1302 1015 1303
rect 488 1203 490 1207
rect 490 1203 493 1207
rect 498 1203 501 1207
rect 501 1203 503 1207
rect 488 1202 493 1203
rect 498 1202 503 1203
rect 1000 1103 1002 1107
rect 1002 1103 1005 1107
rect 1010 1103 1013 1107
rect 1013 1103 1015 1107
rect 1000 1102 1005 1103
rect 1010 1102 1015 1103
rect 488 1003 490 1007
rect 490 1003 493 1007
rect 498 1003 501 1007
rect 501 1003 503 1007
rect 488 1002 493 1003
rect 498 1002 503 1003
rect 1000 903 1002 907
rect 1002 903 1005 907
rect 1010 903 1013 907
rect 1013 903 1015 907
rect 1000 902 1005 903
rect 1010 902 1015 903
rect 488 803 490 807
rect 490 803 493 807
rect 498 803 501 807
rect 501 803 503 807
rect 488 802 493 803
rect 498 802 503 803
rect 1000 703 1002 707
rect 1002 703 1005 707
rect 1010 703 1013 707
rect 1013 703 1015 707
rect 1000 702 1005 703
rect 1010 702 1015 703
rect 488 603 490 607
rect 490 603 493 607
rect 498 603 501 607
rect 501 603 503 607
rect 488 602 493 603
rect 498 602 503 603
rect 1000 503 1002 507
rect 1002 503 1005 507
rect 1010 503 1013 507
rect 1013 503 1015 507
rect 1000 502 1005 503
rect 1010 502 1015 503
rect 488 403 490 407
rect 490 403 493 407
rect 498 403 501 407
rect 501 403 503 407
rect 488 402 493 403
rect 498 402 503 403
rect 1000 303 1002 307
rect 1002 303 1005 307
rect 1010 303 1013 307
rect 1013 303 1015 307
rect 1000 302 1005 303
rect 1010 302 1015 303
rect 488 203 490 207
rect 490 203 493 207
rect 498 203 501 207
rect 501 203 503 207
rect 488 202 493 203
rect 498 202 503 203
rect 1000 103 1002 107
rect 1002 103 1005 107
rect 1010 103 1013 107
rect 1013 103 1015 107
rect 1000 102 1005 103
rect 1010 102 1015 103
rect 488 3 490 7
rect 490 3 493 7
rect 498 3 501 7
rect 501 3 503 7
rect 488 2 493 3
rect 498 2 503 3
<< metal6 >>
rect 488 1207 504 1330
rect 493 1202 498 1207
rect 503 1202 504 1207
rect 488 1007 504 1202
rect 493 1002 498 1007
rect 503 1002 504 1007
rect 488 807 504 1002
rect 493 802 498 807
rect 503 802 504 807
rect 488 607 504 802
rect 493 602 498 607
rect 503 602 504 607
rect 488 407 504 602
rect 493 402 498 407
rect 503 402 504 407
rect 488 207 504 402
rect 493 202 498 207
rect 503 202 504 207
rect 488 7 504 202
rect 493 2 498 7
rect 503 2 504 7
rect 488 -30 504 2
rect 1000 1307 1016 1330
rect 1005 1302 1010 1307
rect 1015 1302 1016 1307
rect 1000 1107 1016 1302
rect 1005 1102 1010 1107
rect 1015 1102 1016 1107
rect 1000 907 1016 1102
rect 1005 902 1010 907
rect 1015 902 1016 907
rect 1000 707 1016 902
rect 1005 702 1010 707
rect 1015 702 1016 707
rect 1000 507 1016 702
rect 1005 502 1010 507
rect 1015 502 1016 507
rect 1000 307 1016 502
rect 1005 302 1010 307
rect 1015 302 1016 307
rect 1000 107 1016 302
rect 1005 102 1010 107
rect 1015 102 1016 107
rect 1000 -30 1016 102
use XOR2X1  XOR2X1_17
timestamp 1696374713
transform 1 0 4 0 -1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_49
timestamp 1696374713
transform 1 0 60 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_52
timestamp 1696374713
transform -1 0 116 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1696374713
transform 1 0 4 0 1 105
box -2 -3 98 103
use INVX1  INVX1_32
timestamp 1696374713
transform 1 0 100 0 1 105
box -2 -3 18 103
use XOR2X1  XOR2X1_13
timestamp 1696374713
transform -1 0 172 0 -1 105
box -2 -3 58 103
use OAI21X1  OAI21X1_51
timestamp 1696374713
transform -1 0 204 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1696374713
transform -1 0 220 0 -1 105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_19
timestamp 1696374713
transform 1 0 116 0 1 105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1696374713
transform 1 0 172 0 1 105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_17
timestamp 1696374713
transform 1 0 220 0 -1 105
box -2 -3 58 103
use OAI21X1  OAI21X1_50
timestamp 1696374713
transform -1 0 308 0 -1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_18
timestamp 1696374713
transform 1 0 268 0 1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_30
timestamp 1696374713
transform -1 0 332 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_30
timestamp 1696374713
transform -1 0 348 0 -1 105
box -2 -3 18 103
use XOR2X1  XOR2X1_12
timestamp 1696374713
transform 1 0 348 0 -1 105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1696374713
transform 1 0 404 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1696374713
transform 1 0 324 0 1 105
box -2 -3 98 103
use FILL  FILL_0_0_0
timestamp 1696374713
transform 1 0 500 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1696374713
transform 1 0 508 0 -1 105
box -2 -3 10 103
use AND2X2  AND2X2_6
timestamp 1696374713
transform -1 0 452 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_45
timestamp 1696374713
transform -1 0 476 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_46
timestamp 1696374713
transform 1 0 476 0 1 105
box -2 -3 26 103
use FILL  FILL_1_0_0
timestamp 1696374713
transform 1 0 500 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1696374713
transform 1 0 508 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1696374713
transform 1 0 516 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1696374713
transform 1 0 516 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_1
timestamp 1696374713
transform -1 0 636 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1696374713
transform -1 0 732 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1696374713
transform 1 0 612 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_2
timestamp 1696374713
transform 1 0 708 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1696374713
transform -1 0 756 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1696374713
transform -1 0 852 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_1
timestamp 1696374713
transform -1 0 756 0 1 105
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1696374713
transform 1 0 756 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_60
timestamp 1696374713
transform 1 0 772 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_3
timestamp 1696374713
transform -1 0 828 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1696374713
transform 1 0 852 0 -1 105
box -2 -3 98 103
use AND2X2  AND2X2_9
timestamp 1696374713
transform -1 0 860 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_10
timestamp 1696374713
transform -1 0 892 0 1 105
box -2 -3 34 103
use INVX1  INVX1_50
timestamp 1696374713
transform -1 0 908 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_56
timestamp 1696374713
transform -1 0 940 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1696374713
transform 1 0 948 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_1_0
timestamp 1696374713
transform 1 0 972 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1696374713
transform 1 0 980 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1696374713
transform 1 0 988 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_4
timestamp 1696374713
transform 1 0 940 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1696374713
transform 1 0 972 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1696374713
transform -1 0 1004 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1696374713
transform -1 0 1012 0 1 105
box -2 -3 10 103
use INVX1  INVX1_20
timestamp 1696374713
transform -1 0 1028 0 1 105
box -2 -3 18 103
use BUFX2  BUFX2_4
timestamp 1696374713
transform 1 0 1084 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1696374713
transform 1 0 1108 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_70
timestamp 1696374713
transform -1 0 1060 0 1 105
box -2 -3 34 103
use INVX1  INVX1_21
timestamp 1696374713
transform -1 0 1076 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_61
timestamp 1696374713
transform -1 0 1108 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_11
timestamp 1696374713
transform 1 0 1108 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_5
timestamp 1696374713
transform 1 0 1204 0 -1 105
box -2 -3 26 103
use NOR3X1  NOR3X1_1
timestamp 1696374713
transform 1 0 1140 0 1 105
box -2 -3 66 103
use AOI21X1  AOI21X1_57
timestamp 1696374713
transform -1 0 1236 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1696374713
transform 1 0 1228 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_48
timestamp 1696374713
transform 1 0 1236 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_30
timestamp 1696374713
transform 1 0 1260 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_3
timestamp 1696374713
transform -1 0 1348 0 1 105
box -2 -3 58 103
use BUFX2  BUFX2_6
timestamp 1696374713
transform 1 0 1324 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1696374713
transform 1 0 1348 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1696374713
transform 1 0 1348 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_8
timestamp 1696374713
transform 1 0 1444 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1696374713
transform -1 0 1492 0 -1 105
box -2 -3 26 103
use FILL  FILL_1_1
timestamp 1696374713
transform -1 0 1500 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1696374713
transform -1 0 1508 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_3
timestamp 1696374713
transform -1 0 1516 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_7
timestamp 1696374713
transform 1 0 1444 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_46
timestamp 1696374713
transform 1 0 1468 0 1 105
box -2 -3 34 103
use FILL  FILL_2_1
timestamp 1696374713
transform 1 0 1500 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1696374713
transform 1 0 1508 0 1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_5
timestamp 1696374713
transform 1 0 4 0 -1 305
box -2 -3 74 103
use XNOR2X1  XNOR2X1_23
timestamp 1696374713
transform -1 0 132 0 -1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1696374713
transform 1 0 132 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1696374713
transform 1 0 228 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1696374713
transform 1 0 324 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1696374713
transform 1 0 420 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1696374713
transform 1 0 516 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1696374713
transform 1 0 524 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1696374713
transform 1 0 532 0 -1 305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_1
timestamp 1696374713
transform -1 0 700 0 -1 305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_3
timestamp 1696374713
transform 1 0 700 0 -1 305
box -2 -3 74 103
use XNOR2X1  XNOR2X1_1
timestamp 1696374713
transform 1 0 772 0 -1 305
box -2 -3 58 103
use INVX1  INVX1_3
timestamp 1696374713
transform -1 0 844 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_1
timestamp 1696374713
transform -1 0 876 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1696374713
transform -1 0 900 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1696374713
transform 1 0 900 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_6
timestamp 1696374713
transform -1 0 948 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_2
timestamp 1696374713
transform -1 0 980 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1696374713
transform -1 0 1012 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1696374713
transform -1 0 1020 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1696374713
transform -1 0 1028 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_4
timestamp 1696374713
transform -1 0 1060 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_3
timestamp 1696374713
transform -1 0 1092 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_5
timestamp 1696374713
transform -1 0 1108 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_8
timestamp 1696374713
transform 1 0 1108 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_1
timestamp 1696374713
transform 1 0 1132 0 -1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_2
timestamp 1696374713
transform -1 0 1228 0 -1 305
box -2 -3 66 103
use OAI21X1  OAI21X1_21
timestamp 1696374713
transform 1 0 1228 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1696374713
transform 1 0 1260 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_6
timestamp 1696374713
transform 1 0 1284 0 -1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_15
timestamp 1696374713
transform -1 0 1348 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_53
timestamp 1696374713
transform -1 0 1380 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1696374713
transform 1 0 1380 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1696374713
transform -1 0 1436 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_69
timestamp 1696374713
transform 1 0 1436 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_42
timestamp 1696374713
transform -1 0 1500 0 -1 305
box -2 -3 34 103
use FILL  FILL_3_1
timestamp 1696374713
transform -1 0 1508 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1696374713
transform -1 0 1516 0 -1 305
box -2 -3 10 103
use XOR2X1  XOR2X1_15
timestamp 1696374713
transform 1 0 4 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_53
timestamp 1696374713
transform 1 0 60 0 1 305
box -2 -3 26 103
use INVX1  INVX1_38
timestamp 1696374713
transform -1 0 100 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_55
timestamp 1696374713
transform -1 0 132 0 1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_16
timestamp 1696374713
transform -1 0 188 0 1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1696374713
transform 1 0 188 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1696374713
transform 1 0 284 0 1 305
box -2 -3 98 103
use INVX1  INVX1_40
timestamp 1696374713
transform -1 0 396 0 1 305
box -2 -3 18 103
use XOR2X1  XOR2X1_18
timestamp 1696374713
transform -1 0 452 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_54
timestamp 1696374713
transform -1 0 476 0 1 305
box -2 -3 26 103
use FILL  FILL_3_0_0
timestamp 1696374713
transform 1 0 476 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1696374713
transform 1 0 484 0 1 305
box -2 -3 10 103
use XOR2X1  XOR2X1_19
timestamp 1696374713
transform 1 0 492 0 1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1696374713
transform 1 0 548 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1696374713
transform 1 0 644 0 1 305
box -2 -3 98 103
use INVX4  INVX4_1
timestamp 1696374713
transform 1 0 740 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_19
timestamp 1696374713
transform -1 0 788 0 1 305
box -2 -3 26 103
use INVX1  INVX1_11
timestamp 1696374713
transform 1 0 788 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_2
timestamp 1696374713
transform 1 0 804 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_4
timestamp 1696374713
transform -1 0 860 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_59
timestamp 1696374713
transform -1 0 892 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1
timestamp 1696374713
transform -1 0 924 0 1 305
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1696374713
transform -1 0 940 0 1 305
box -2 -3 18 103
use BUFX4  BUFX4_1
timestamp 1696374713
transform 1 0 940 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1696374713
transform 1 0 972 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1696374713
transform -1 0 1012 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1696374713
transform -1 0 1020 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_8
timestamp 1696374713
transform -1 0 1044 0 1 305
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1696374713
transform 1 0 1044 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_3
timestamp 1696374713
transform -1 0 1092 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1696374713
transform 1 0 1092 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_14
timestamp 1696374713
transform 1 0 1124 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_10
timestamp 1696374713
transform -1 0 1188 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1696374713
transform -1 0 1212 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_45
timestamp 1696374713
transform 1 0 1212 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1696374713
transform -1 0 1276 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_71
timestamp 1696374713
transform -1 0 1308 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_27
timestamp 1696374713
transform 1 0 1308 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_32
timestamp 1696374713
transform -1 0 1372 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_72
timestamp 1696374713
transform -1 0 1404 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_49
timestamp 1696374713
transform 1 0 1404 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_74
timestamp 1696374713
transform 1 0 1436 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_44
timestamp 1696374713
transform -1 0 1500 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1696374713
transform 1 0 1500 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1696374713
transform 1 0 1508 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_48
timestamp 1696374713
transform 1 0 4 0 -1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_14
timestamp 1696374713
transform -1 0 84 0 -1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_49
timestamp 1696374713
transform -1 0 116 0 -1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_11
timestamp 1696374713
transform -1 0 172 0 -1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1696374713
transform 1 0 172 0 -1 505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_2
timestamp 1696374713
transform -1 0 340 0 -1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_33
timestamp 1696374713
transform -1 0 364 0 -1 505
box -2 -3 26 103
use AND2X2  AND2X2_7
timestamp 1696374713
transform 1 0 364 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_56
timestamp 1696374713
transform 1 0 396 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1696374713
transform -1 0 444 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_34
timestamp 1696374713
transform 1 0 444 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_54
timestamp 1696374713
transform -1 0 500 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_0_0
timestamp 1696374713
transform -1 0 508 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1696374713
transform -1 0 516 0 -1 505
box -2 -3 10 103
use XOR2X1  XOR2X1_20
timestamp 1696374713
transform -1 0 572 0 -1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1696374713
transform 1 0 572 0 -1 505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_4
timestamp 1696374713
transform -1 0 740 0 -1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_9
timestamp 1696374713
transform 1 0 740 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_7
timestamp 1696374713
transform -1 0 796 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1696374713
transform -1 0 812 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_8
timestamp 1696374713
transform -1 0 844 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_1
timestamp 1696374713
transform 1 0 844 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_10
timestamp 1696374713
transform 1 0 860 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_16
timestamp 1696374713
transform 1 0 884 0 -1 505
box -2 -3 26 103
use BUFX4  BUFX4_3
timestamp 1696374713
transform 1 0 908 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1696374713
transform 1 0 940 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_5
timestamp 1696374713
transform -1 0 988 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1696374713
transform -1 0 1012 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_1_0
timestamp 1696374713
transform -1 0 1020 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1696374713
transform -1 0 1028 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_7
timestamp 1696374713
transform -1 0 1060 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_9
timestamp 1696374713
transform -1 0 1076 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_3
timestamp 1696374713
transform 1 0 1076 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1696374713
transform 1 0 1108 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1696374713
transform 1 0 1140 0 -1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_16
timestamp 1696374713
transform -1 0 1188 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1696374713
transform 1 0 1188 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_5
timestamp 1696374713
transform 1 0 1220 0 -1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_20
timestamp 1696374713
transform 1 0 1236 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1696374713
transform 1 0 1268 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1696374713
transform -1 0 1332 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_21
timestamp 1696374713
transform -1 0 1364 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1696374713
transform 1 0 1364 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1696374713
transform 1 0 1396 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_73
timestamp 1696374713
transform 1 0 1420 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1696374713
transform 1 0 1452 0 -1 505
box -2 -3 26 103
use AND2X2  AND2X2_1
timestamp 1696374713
transform 1 0 1476 0 -1 505
box -2 -3 34 103
use FILL  FILL_5_1
timestamp 1696374713
transform -1 0 1516 0 -1 505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_16
timestamp 1696374713
transform 1 0 4 0 1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1696374713
transform 1 0 60 0 1 505
box -2 -3 98 103
use XNOR2X1  XNOR2X1_26
timestamp 1696374713
transform 1 0 156 0 1 505
box -2 -3 58 103
use NAND2X1  NAND2X1_59
timestamp 1696374713
transform 1 0 212 0 1 505
box -2 -3 26 103
use INVX1  INVX1_47
timestamp 1696374713
transform 1 0 236 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_42
timestamp 1696374713
transform 1 0 252 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_43
timestamp 1696374713
transform 1 0 276 0 1 505
box -2 -3 26 103
use INVX1  INVX1_48
timestamp 1696374713
transform 1 0 300 0 1 505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_6
timestamp 1696374713
transform -1 0 388 0 1 505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1696374713
transform 1 0 388 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1696374713
transform 1 0 484 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1696374713
transform 1 0 492 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_12
timestamp 1696374713
transform 1 0 500 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_8
timestamp 1696374713
transform -1 0 564 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_9
timestamp 1696374713
transform 1 0 564 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_15
timestamp 1696374713
transform 1 0 588 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_10
timestamp 1696374713
transform 1 0 612 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_5
timestamp 1696374713
transform -1 0 660 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_6
timestamp 1696374713
transform 1 0 660 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_22
timestamp 1696374713
transform 1 0 692 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1696374713
transform 1 0 724 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1696374713
transform -1 0 772 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_4
timestamp 1696374713
transform 1 0 772 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_3
timestamp 1696374713
transform -1 0 820 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_5
timestamp 1696374713
transform 1 0 820 0 1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1696374713
transform 1 0 844 0 1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_9
timestamp 1696374713
transform -1 0 916 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1696374713
transform 1 0 916 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1696374713
transform -1 0 980 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_8
timestamp 1696374713
transform 1 0 980 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1696374713
transform 1 0 1012 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1696374713
transform 1 0 1020 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_15
timestamp 1696374713
transform 1 0 1028 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_29
timestamp 1696374713
transform -1 0 1092 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_17
timestamp 1696374713
transform 1 0 1092 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1696374713
transform 1 0 1124 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_28
timestamp 1696374713
transform -1 0 1188 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_19
timestamp 1696374713
transform 1 0 1188 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_22
timestamp 1696374713
transform -1 0 1252 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_18
timestamp 1696374713
transform -1 0 1284 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_32
timestamp 1696374713
transform 1 0 1284 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_52
timestamp 1696374713
transform -1 0 1348 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_50
timestamp 1696374713
transform 1 0 1348 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1696374713
transform 1 0 1380 0 1 505
box -2 -3 26 103
use INVX2  INVX2_7
timestamp 1696374713
transform -1 0 1420 0 1 505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_12
timestamp 1696374713
transform -1 0 1476 0 1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_33
timestamp 1696374713
transform 1 0 1476 0 1 505
box -2 -3 34 103
use FILL  FILL_6_1
timestamp 1696374713
transform 1 0 1508 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_26
timestamp 1696374713
transform 1 0 4 0 -1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_15
timestamp 1696374713
transform -1 0 84 0 -1 705
box -2 -3 58 103
use INVX1  INVX1_29
timestamp 1696374713
transform 1 0 84 0 -1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_51
timestamp 1696374713
transform 1 0 100 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1696374713
transform -1 0 156 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_50
timestamp 1696374713
transform -1 0 180 0 -1 705
box -2 -3 26 103
use XOR2X1  XOR2X1_14
timestamp 1696374713
transform -1 0 236 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_10
timestamp 1696374713
transform -1 0 292 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_22
timestamp 1696374713
transform -1 0 348 0 -1 705
box -2 -3 58 103
use NOR2X1  NOR2X1_44
timestamp 1696374713
transform 1 0 348 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1696374713
transform 1 0 372 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_0_0
timestamp 1696374713
transform 1 0 468 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1696374713
transform 1 0 476 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1696374713
transform 1 0 484 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_33
timestamp 1696374713
transform 1 0 580 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_16
timestamp 1696374713
transform 1 0 604 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_18
timestamp 1696374713
transform -1 0 660 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1696374713
transform -1 0 692 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1696374713
transform 1 0 692 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_19
timestamp 1696374713
transform -1 0 740 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_16
timestamp 1696374713
transform 1 0 740 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1696374713
transform 1 0 772 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_18
timestamp 1696374713
transform 1 0 796 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_2
timestamp 1696374713
transform -1 0 852 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_4
timestamp 1696374713
transform 1 0 852 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1696374713
transform -1 0 908 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_2
timestamp 1696374713
transform 1 0 908 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_11
timestamp 1696374713
transform -1 0 980 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_9
timestamp 1696374713
transform 1 0 980 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1696374713
transform 1 0 1012 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1696374713
transform 1 0 1020 0 -1 705
box -2 -3 10 103
use INVX2  INVX2_3
timestamp 1696374713
transform 1 0 1028 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_10
timestamp 1696374713
transform -1 0 1076 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_12
timestamp 1696374713
transform 1 0 1076 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1696374713
transform 1 0 1108 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_24
timestamp 1696374713
transform 1 0 1140 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1696374713
transform -1 0 1204 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_20
timestamp 1696374713
transform 1 0 1204 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1696374713
transform 1 0 1236 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1696374713
transform 1 0 1268 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1696374713
transform 1 0 1300 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1696374713
transform 1 0 1332 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1696374713
transform 1 0 1364 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_48
timestamp 1696374713
transform -1 0 1428 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_51
timestamp 1696374713
transform -1 0 1460 0 -1 705
box -2 -3 34 103
use XOR2X1  XOR2X1_1
timestamp 1696374713
transform -1 0 1516 0 -1 705
box -2 -3 58 103
use INVX1  INVX1_27
timestamp 1696374713
transform 1 0 4 0 1 705
box -2 -3 18 103
use INVX1  INVX1_28
timestamp 1696374713
transform 1 0 20 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_25
timestamp 1696374713
transform 1 0 36 0 1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_20
timestamp 1696374713
transform 1 0 60 0 1 705
box -2 -3 58 103
use INVX1  INVX1_33
timestamp 1696374713
transform 1 0 116 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_53
timestamp 1696374713
transform 1 0 132 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_53
timestamp 1696374713
transform -1 0 196 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1696374713
transform 1 0 196 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1696374713
transform 1 0 292 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1696374713
transform 1 0 388 0 1 705
box -2 -3 98 103
use FILL  FILL_7_0_0
timestamp 1696374713
transform 1 0 484 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1696374713
transform 1 0 492 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1696374713
transform 1 0 500 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_17
timestamp 1696374713
transform 1 0 596 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_9
timestamp 1696374713
transform -1 0 652 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_11
timestamp 1696374713
transform -1 0 684 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1696374713
transform 1 0 684 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_24
timestamp 1696374713
transform -1 0 740 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1696374713
transform 1 0 740 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1696374713
transform 1 0 772 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1696374713
transform 1 0 804 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1696374713
transform 1 0 836 0 1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_1
timestamp 1696374713
transform 1 0 860 0 1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_11
timestamp 1696374713
transform 1 0 900 0 1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_2
timestamp 1696374713
transform -1 0 964 0 1 705
box -2 -3 42 103
use AOI21X1  AOI21X1_6
timestamp 1696374713
transform 1 0 964 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1696374713
transform 1 0 996 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1696374713
transform 1 0 1004 0 1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_5
timestamp 1696374713
transform 1 0 1012 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1696374713
transform 1 0 1044 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_7
timestamp 1696374713
transform 1 0 1068 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_22
timestamp 1696374713
transform 1 0 1092 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_13
timestamp 1696374713
transform -1 0 1148 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1696374713
transform -1 0 1180 0 1 705
box -2 -3 34 103
use INVX2  INVX2_4
timestamp 1696374713
transform -1 0 1196 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_19
timestamp 1696374713
transform 1 0 1196 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_22
timestamp 1696374713
transform 1 0 1228 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1696374713
transform 1 0 1260 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_23
timestamp 1696374713
transform 1 0 1292 0 1 705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1696374713
transform 1 0 1324 0 1 705
box -2 -3 58 103
use NAND3X1  NAND3X1_49
timestamp 1696374713
transform 1 0 1380 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_47
timestamp 1696374713
transform 1 0 1412 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_44
timestamp 1696374713
transform -1 0 1476 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_44
timestamp 1696374713
transform 1 0 1476 0 1 705
box -2 -3 34 103
use FILL  FILL_8_1
timestamp 1696374713
transform 1 0 1508 0 1 705
box -2 -3 10 103
use INVX1  INVX1_36
timestamp 1696374713
transform 1 0 4 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_52
timestamp 1696374713
transform 1 0 20 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1696374713
transform 1 0 44 0 -1 905
box -2 -3 34 103
use AND2X2  AND2X2_5
timestamp 1696374713
transform 1 0 76 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_54
timestamp 1696374713
transform -1 0 140 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1696374713
transform 1 0 140 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_52
timestamp 1696374713
transform -1 0 188 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1696374713
transform 1 0 188 0 -1 905
box -2 -3 26 103
use INVX2  INVX2_8
timestamp 1696374713
transform 1 0 212 0 -1 905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_21
timestamp 1696374713
transform -1 0 284 0 -1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1696374713
transform 1 0 284 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1696374713
transform 1 0 380 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_0_0
timestamp 1696374713
transform 1 0 476 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1696374713
transform 1 0 484 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1696374713
transform 1 0 492 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_49
timestamp 1696374713
transform 1 0 588 0 -1 905
box -2 -3 18 103
use AND2X2  AND2X2_8
timestamp 1696374713
transform 1 0 604 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1696374713
transform 1 0 636 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_34
timestamp 1696374713
transform 1 0 660 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_27
timestamp 1696374713
transform -1 0 708 0 -1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_3
timestamp 1696374713
transform -1 0 748 0 -1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_35
timestamp 1696374713
transform 1 0 748 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_26
timestamp 1696374713
transform 1 0 772 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1696374713
transform -1 0 828 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1696374713
transform -1 0 844 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_35
timestamp 1696374713
transform 1 0 844 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_19
timestamp 1696374713
transform 1 0 876 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_15
timestamp 1696374713
transform 1 0 900 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_27
timestamp 1696374713
transform 1 0 916 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1696374713
transform -1 0 988 0 -1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_20
timestamp 1696374713
transform 1 0 988 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_1_0
timestamp 1696374713
transform -1 0 1020 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1696374713
transform -1 0 1028 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_21
timestamp 1696374713
transform -1 0 1052 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_12
timestamp 1696374713
transform 1 0 1052 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1696374713
transform 1 0 1084 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1696374713
transform 1 0 1116 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1696374713
transform 1 0 1148 0 -1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_3
timestamp 1696374713
transform 1 0 1180 0 -1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_12
timestamp 1696374713
transform 1 0 1220 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_18
timestamp 1696374713
transform -1 0 1276 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1696374713
transform 1 0 1276 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1696374713
transform -1 0 1340 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_46
timestamp 1696374713
transform -1 0 1372 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_43
timestamp 1696374713
transform -1 0 1404 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_30
timestamp 1696374713
transform 1 0 1404 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_45
timestamp 1696374713
transform 1 0 1436 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_40
timestamp 1696374713
transform 1 0 1468 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1696374713
transform -1 0 1508 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1696374713
transform -1 0 1516 0 -1 905
box -2 -3 10 103
use INVX1  INVX1_34
timestamp 1696374713
transform 1 0 4 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_51
timestamp 1696374713
transform -1 0 44 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_31
timestamp 1696374713
transform 1 0 44 0 1 905
box -2 -3 26 103
use INVX1  INVX1_35
timestamp 1696374713
transform 1 0 68 0 1 905
box -2 -3 18 103
use AND2X2  AND2X2_4
timestamp 1696374713
transform 1 0 84 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_22
timestamp 1696374713
transform -1 0 172 0 1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1696374713
transform 1 0 172 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1696374713
transform 1 0 268 0 1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_38
timestamp 1696374713
transform 1 0 364 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_57
timestamp 1696374713
transform 1 0 388 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1696374713
transform 1 0 412 0 1 905
box -2 -3 98 103
use FILL  FILL_9_0_0
timestamp 1696374713
transform 1 0 508 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1696374713
transform 1 0 516 0 1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_39
timestamp 1696374713
transform 1 0 524 0 1 905
box -2 -3 26 103
use INVX1  INVX1_45
timestamp 1696374713
transform -1 0 564 0 1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_55
timestamp 1696374713
transform -1 0 596 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_75
timestamp 1696374713
transform 1 0 596 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_11
timestamp 1696374713
transform 1 0 628 0 1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_4
timestamp 1696374713
transform 1 0 652 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_31
timestamp 1696374713
transform 1 0 692 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_25
timestamp 1696374713
transform 1 0 724 0 1 905
box -2 -3 34 103
use INVX1  INVX1_12
timestamp 1696374713
transform -1 0 772 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_24
timestamp 1696374713
transform -1 0 804 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1696374713
transform 1 0 804 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1696374713
transform 1 0 836 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_32
timestamp 1696374713
transform 1 0 860 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_38
timestamp 1696374713
transform -1 0 908 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_54
timestamp 1696374713
transform 1 0 908 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_36
timestamp 1696374713
transform 1 0 940 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_31
timestamp 1696374713
transform 1 0 964 0 1 905
box -2 -3 26 103
use FILL  FILL_9_1_0
timestamp 1696374713
transform 1 0 988 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1696374713
transform 1 0 996 0 1 905
box -2 -3 10 103
use OAI22X1  OAI22X1_5
timestamp 1696374713
transform 1 0 1004 0 1 905
box -2 -3 42 103
use AOI22X1  AOI22X1_5
timestamp 1696374713
transform 1 0 1044 0 1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_29
timestamp 1696374713
transform 1 0 1084 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_31
timestamp 1696374713
transform 1 0 1108 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_26
timestamp 1696374713
transform 1 0 1140 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1696374713
transform -1 0 1196 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_29
timestamp 1696374713
transform 1 0 1196 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_38
timestamp 1696374713
transform 1 0 1228 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_35
timestamp 1696374713
transform -1 0 1292 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_42
timestamp 1696374713
transform -1 0 1324 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_39
timestamp 1696374713
transform -1 0 1356 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_41
timestamp 1696374713
transform 1 0 1356 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_36
timestamp 1696374713
transform 1 0 1388 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1696374713
transform 1 0 1420 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1696374713
transform 1 0 1452 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_68
timestamp 1696374713
transform -1 0 1508 0 1 905
box -2 -3 34 103
use FILL  FILL_10_1
timestamp 1696374713
transform 1 0 1508 0 1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_23
timestamp 1696374713
transform 1 0 4 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_24
timestamp 1696374713
transform 1 0 28 0 -1 1105
box -2 -3 18 103
use INVX1  INVX1_25
timestamp 1696374713
transform 1 0 44 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_22
timestamp 1696374713
transform -1 0 84 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_47
timestamp 1696374713
transform 1 0 84 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1696374713
transform 1 0 108 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1696374713
transform 1 0 204 0 -1 1105
box -2 -3 98 103
use XOR2X1  XOR2X1_6
timestamp 1696374713
transform 1 0 300 0 -1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_55
timestamp 1696374713
transform 1 0 356 0 -1 1105
box -2 -3 26 103
use XOR2X1  XOR2X1_21
timestamp 1696374713
transform -1 0 436 0 -1 1105
box -2 -3 58 103
use INVX1  INVX1_41
timestamp 1696374713
transform 1 0 436 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_57
timestamp 1696374713
transform -1 0 484 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1696374713
transform -1 0 492 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1696374713
transform -1 0 500 0 -1 1105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_24
timestamp 1696374713
transform -1 0 556 0 -1 1105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1696374713
transform 1 0 556 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1696374713
transform 1 0 652 0 -1 1105
box -2 -3 98 103
use XOR2X1  XOR2X1_3
timestamp 1696374713
transform 1 0 748 0 -1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_37
timestamp 1696374713
transform 1 0 804 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1696374713
transform 1 0 828 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_55
timestamp 1696374713
transform -1 0 892 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_56
timestamp 1696374713
transform -1 0 924 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_37
timestamp 1696374713
transform -1 0 956 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_25
timestamp 1696374713
transform 1 0 956 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1696374713
transform 1 0 988 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1696374713
transform -1 0 1020 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1696374713
transform -1 0 1028 0 -1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_32
timestamp 1696374713
transform -1 0 1060 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_33
timestamp 1696374713
transform -1 0 1092 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1696374713
transform 1 0 1092 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_28
timestamp 1696374713
transform -1 0 1140 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1696374713
transform 1 0 1140 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_34
timestamp 1696374713
transform -1 0 1204 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_42
timestamp 1696374713
transform 1 0 1204 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_40
timestamp 1696374713
transform 1 0 1236 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1696374713
transform -1 0 1300 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1696374713
transform 1 0 1300 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1696374713
transform -1 0 1364 0 -1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_4
timestamp 1696374713
transform -1 0 1420 0 -1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_41
timestamp 1696374713
transform 1 0 1420 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_67
timestamp 1696374713
transform -1 0 1484 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_47
timestamp 1696374713
transform 1 0 1484 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_45
timestamp 1696374713
transform 1 0 4 0 1 1105
box -2 -3 26 103
use XOR2X1  XOR2X1_8
timestamp 1696374713
transform -1 0 84 0 1 1105
box -2 -3 58 103
use NOR2X1  NOR2X1_24
timestamp 1696374713
transform 1 0 84 0 1 1105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_13
timestamp 1696374713
transform -1 0 164 0 1 1105
box -2 -3 58 103
use INVX1  INVX1_26
timestamp 1696374713
transform 1 0 164 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_48
timestamp 1696374713
transform 1 0 180 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1696374713
transform -1 0 236 0 1 1105
box -2 -3 26 103
use XOR2X1  XOR2X1_9
timestamp 1696374713
transform -1 0 292 0 1 1105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1696374713
transform 1 0 292 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_36
timestamp 1696374713
transform -1 0 412 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_42
timestamp 1696374713
transform 1 0 412 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_43
timestamp 1696374713
transform 1 0 428 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_37
timestamp 1696374713
transform 1 0 444 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_35
timestamp 1696374713
transform 1 0 468 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_0_0
timestamp 1696374713
transform 1 0 492 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1696374713
transform 1 0 500 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_58
timestamp 1696374713
transform 1 0 508 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_58
timestamp 1696374713
transform 1 0 540 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_40
timestamp 1696374713
transform 1 0 564 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_41
timestamp 1696374713
transform 1 0 588 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_46
timestamp 1696374713
transform -1 0 628 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1696374713
transform 1 0 628 0 1 1105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_5
timestamp 1696374713
transform 1 0 724 0 1 1105
box -2 -3 58 103
use NOR3X1  NOR3X1_3
timestamp 1696374713
transform -1 0 844 0 1 1105
box -2 -3 66 103
use OAI21X1  OAI21X1_35
timestamp 1696374713
transform 1 0 844 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_17
timestamp 1696374713
transform -1 0 892 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_59
timestamp 1696374713
transform 1 0 892 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1696374713
transform 1 0 924 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_57
timestamp 1696374713
transform -1 0 972 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_41
timestamp 1696374713
transform -1 0 1004 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_1_0
timestamp 1696374713
transform 1 0 1004 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1696374713
transform 1 0 1012 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_36
timestamp 1696374713
transform 1 0 1020 0 1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_5
timestamp 1696374713
transform 1 0 1052 0 1 1105
box -2 -3 66 103
use OAI21X1  OAI21X1_39
timestamp 1696374713
transform 1 0 1116 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_10
timestamp 1696374713
transform 1 0 1148 0 1 1105
box -2 -3 58 103
use NAND3X1  NAND3X1_64
timestamp 1696374713
transform 1 0 1204 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1696374713
transform -1 0 1268 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_43
timestamp 1696374713
transform 1 0 1268 0 1 1105
box -2 -3 34 103
use XOR2X1  XOR2X1_2
timestamp 1696374713
transform -1 0 1356 0 1 1105
box -2 -3 58 103
use NAND3X1  NAND3X1_62
timestamp 1696374713
transform -1 0 1388 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1696374713
transform 1 0 1388 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_63
timestamp 1696374713
transform -1 0 1452 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1696374713
transform -1 0 1468 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_33
timestamp 1696374713
transform -1 0 1500 0 1 1105
box -2 -3 34 103
use FILL  FILL_12_1
timestamp 1696374713
transform 1 0 1500 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1696374713
transform 1 0 1508 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_20
timestamp 1696374713
transform -1 0 28 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1696374713
transform 1 0 28 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1696374713
transform 1 0 60 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_50
timestamp 1696374713
transform -1 0 116 0 -1 1305
box -2 -3 34 103
use XOR2X1  XOR2X1_7
timestamp 1696374713
transform -1 0 172 0 -1 1305
box -2 -3 58 103
use OAI21X1  OAI21X1_47
timestamp 1696374713
transform -1 0 204 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_23
timestamp 1696374713
transform -1 0 220 0 -1 1305
box -2 -3 18 103
use INVX1  INVX1_22
timestamp 1696374713
transform -1 0 236 0 -1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_5
timestamp 1696374713
transform -1 0 292 0 -1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_44
timestamp 1696374713
transform -1 0 316 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1696374713
transform 1 0 316 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_29
timestamp 1696374713
transform -1 0 436 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1696374713
transform -1 0 468 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_28
timestamp 1696374713
transform -1 0 492 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_0_0
timestamp 1696374713
transform 1 0 492 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1696374713
transform 1 0 500 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_56
timestamp 1696374713
transform 1 0 508 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_44
timestamp 1696374713
transform 1 0 532 0 -1 1305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_25
timestamp 1696374713
transform -1 0 604 0 -1 1305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1696374713
transform 1 0 604 0 -1 1305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_7
timestamp 1696374713
transform -1 0 756 0 -1 1305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_6
timestamp 1696374713
transform 1 0 756 0 -1 1305
box -2 -3 58 103
use INVX2  INVX2_6
timestamp 1696374713
transform 1 0 812 0 -1 1305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_8
timestamp 1696374713
transform -1 0 884 0 -1 1305
box -2 -3 58 103
use NAND3X1  NAND3X1_60
timestamp 1696374713
transform 1 0 884 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_38
timestamp 1696374713
transform -1 0 948 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1696374713
transform -1 0 980 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_37
timestamp 1696374713
transform -1 0 1012 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_1_0
timestamp 1696374713
transform -1 0 1020 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1696374713
transform -1 0 1028 0 -1 1305
box -2 -3 10 103
use NOR3X1  NOR3X1_4
timestamp 1696374713
transform -1 0 1092 0 -1 1305
box -2 -3 66 103
use OAI21X1  OAI21X1_36
timestamp 1696374713
transform 1 0 1092 0 -1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_9
timestamp 1696374713
transform -1 0 1180 0 -1 1305
box -2 -3 58 103
use AOI21X1  AOI21X1_46
timestamp 1696374713
transform 1 0 1180 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1696374713
transform 1 0 1212 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_66
timestamp 1696374713
transform 1 0 1228 0 -1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_11
timestamp 1696374713
transform -1 0 1316 0 -1 1305
box -2 -3 58 103
use NAND3X1  NAND3X1_65
timestamp 1696374713
transform 1 0 1316 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_45
timestamp 1696374713
transform -1 0 1380 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1696374713
transform 1 0 1380 0 -1 1305
box -2 -3 34 103
use XOR2X1  XOR2X1_4
timestamp 1696374713
transform -1 0 1468 0 -1 1305
box -2 -3 58 103
use NOR2X1  NOR2X1_17
timestamp 1696374713
transform 1 0 1468 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1696374713
transform -1 0 1500 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1696374713
transform -1 0 1508 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_3
timestamp 1696374713
transform -1 0 1516 0 -1 1305
box -2 -3 10 103
<< labels >>
flabel metal6 s 488 -30 504 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1000 -30 1016 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 454 1328 458 1332 3 FreeSans 24 90 0 0 A[0]
port 2 nsew
flabel metal2 s 214 1328 218 1332 3 FreeSans 24 90 0 0 A[1]
port 3 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 90 0 0 A[2]
port 4 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 A[3]
port 5 nsew
flabel metal3 s -26 1168 -22 1172 7 FreeSans 24 0 0 0 A[4]
port 6 nsew
flabel metal3 s -26 658 -22 662 7 FreeSans 24 0 0 0 A[5]
port 7 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 A[6]
port 8 nsew
flabel metal3 s -26 678 -22 682 7 FreeSans 24 0 0 0 A[7]
port 9 nsew
flabel metal2 s 478 1328 482 1332 3 FreeSans 24 90 0 0 B[0]
port 10 nsew
flabel metal2 s 238 1328 242 1332 3 FreeSans 24 90 0 0 B[1]
port 11 nsew
flabel metal3 s -26 1268 -22 1272 7 FreeSans 24 90 0 0 B[2]
port 12 nsew
flabel metal3 s -26 1068 -22 1072 7 FreeSans 24 0 0 0 B[3]
port 13 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 B[4]
port 14 nsew
flabel metal3 s -26 778 -22 782 7 FreeSans 24 0 0 0 B[5]
port 15 nsew
flabel metal3 s -26 468 -22 472 7 FreeSans 24 0 0 0 B[6]
port 16 nsew
flabel metal3 s -26 698 -22 702 7 FreeSans 24 0 0 0 B[7]
port 17 nsew
flabel metal2 s 358 -22 362 -18 7 FreeSans 24 270 0 0 C[0]
port 18 nsew
flabel metal2 s 238 -22 242 -18 7 FreeSans 24 270 0 0 C[1]
port 19 nsew
flabel metal3 s -26 128 -22 132 7 FreeSans 24 0 0 0 C[2]
port 20 nsew
flabel metal3 s -26 738 -22 742 7 FreeSans 24 0 0 0 C[3]
port 21 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 C[4]
port 22 nsew
flabel metal3 s -26 868 -22 872 7 FreeSans 24 0 0 0 C[5]
port 23 nsew
flabel metal3 s -26 358 -22 362 7 FreeSans 24 0 0 0 C[6]
port 24 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 C[7]
port 25 nsew
flabel metal2 s 430 -22 434 -18 7 FreeSans 24 270 0 0 D[0]
port 26 nsew
flabel metal2 s 542 -22 546 -18 7 FreeSans 24 270 0 0 D[1]
port 27 nsew
flabel metal2 s 102 -22 106 -18 7 FreeSans 24 270 0 0 D[2]
port 28 nsew
flabel metal3 s -26 758 -22 762 7 FreeSans 24 0 0 0 D[3]
port 29 nsew
flabel metal3 s -26 968 -22 972 7 FreeSans 24 0 0 0 D[4]
port 30 nsew
flabel metal3 s -26 848 -22 852 7 FreeSans 24 0 0 0 D[5]
port 31 nsew
flabel metal3 s -26 338 -22 342 7 FreeSans 24 0 0 0 D[6]
port 32 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 D[7]
port 33 nsew
flabel metal3 s -26 268 -22 272 7 FreeSans 24 0 0 0 clk
port 34 nsew
flabel metal2 s 622 -22 626 -18 7 FreeSans 24 270 0 0 F[0]
port 35 nsew
flabel metal2 s 742 -22 746 -18 7 FreeSans 24 270 0 0 F[1]
port 36 nsew
flabel metal2 s 958 -22 962 -18 7 FreeSans 24 270 0 0 F[2]
port 37 nsew
flabel metal2 s 1094 -22 1098 -18 7 FreeSans 24 270 0 0 F[3]
port 38 nsew
flabel metal2 s 1214 -22 1218 -18 7 FreeSans 24 270 0 0 F[4]
port 39 nsew
flabel metal2 s 1334 -22 1338 -18 7 FreeSans 24 270 0 0 F[5]
port 40 nsew
flabel metal3 s 1542 148 1546 152 3 FreeSans 24 0 0 0 F[6]
port 41 nsew
flabel metal2 s 1454 -22 1458 -18 3 FreeSans 24 270 0 0 F[7]
port 42 nsew
<< end >>
