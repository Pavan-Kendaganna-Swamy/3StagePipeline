VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipeline
  CLASS BLOCK ;
  FOREIGN pipeline ;
  ORIGIN 2.600 3.000 ;
  SIZE 157.200 BY 136.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 2.200 120.800 2.600 125.100 ;
        RECT 3.000 120.800 3.400 123.100 ;
        RECT 4.600 120.800 5.000 124.900 ;
        RECT 6.200 120.800 6.600 125.100 ;
        RECT 10.200 120.800 10.600 124.500 ;
        RECT 12.600 120.800 13.100 124.400 ;
        RECT 15.700 121.100 16.200 124.400 ;
        RECT 15.700 120.800 16.100 121.100 ;
        RECT 17.700 120.800 18.100 123.100 ;
        RECT 19.800 120.800 20.200 125.100 ;
        RECT 21.400 120.800 21.800 123.100 ;
        RECT 23.000 120.800 23.400 123.100 ;
        RECT 24.600 120.800 25.100 124.400 ;
        RECT 27.700 121.100 28.200 124.400 ;
        RECT 27.700 120.800 28.100 121.100 ;
        RECT 29.400 120.800 29.800 123.100 ;
        RECT 31.000 120.800 31.400 123.100 ;
        RECT 32.600 120.800 33.000 125.000 ;
        RECT 35.400 120.800 35.800 123.100 ;
        RECT 37.000 120.800 37.400 123.100 ;
        RECT 39.800 120.800 40.200 125.100 ;
        RECT 43.000 120.800 43.400 125.100 ;
        RECT 44.600 120.800 45.000 124.900 ;
        RECT 46.200 120.800 46.600 123.100 ;
        RECT 48.600 120.800 49.000 125.100 ;
        RECT 51.000 120.800 51.400 123.100 ;
        RECT 52.600 120.800 53.000 123.100 ;
        RECT 53.400 120.800 53.800 123.100 ;
        RECT 55.800 120.800 56.300 124.400 ;
        RECT 58.900 121.100 59.400 124.400 ;
        RECT 58.900 120.800 59.300 121.100 ;
        RECT 61.400 120.800 61.800 125.000 ;
        RECT 64.200 120.800 64.600 123.100 ;
        RECT 65.800 120.800 66.200 123.100 ;
        RECT 68.600 120.800 69.000 125.100 ;
        RECT 71.000 120.800 71.500 124.400 ;
        RECT 74.100 121.100 74.600 124.400 ;
        RECT 76.600 121.100 77.100 124.400 ;
        RECT 74.100 120.800 74.500 121.100 ;
        RECT 76.700 120.800 77.100 121.100 ;
        RECT 79.700 120.800 80.200 124.400 ;
        RECT 81.400 120.800 81.800 125.100 ;
        RECT 83.800 120.800 84.300 124.400 ;
        RECT 86.900 121.100 87.400 124.400 ;
        RECT 86.900 120.800 87.300 121.100 ;
        RECT 88.600 120.800 89.000 123.100 ;
        RECT 90.200 120.800 90.600 122.900 ;
        RECT 92.100 120.800 92.500 123.100 ;
        RECT 94.200 120.800 94.600 125.100 ;
        RECT 95.800 120.800 96.200 122.900 ;
        RECT 97.400 120.800 97.800 123.100 ;
        RECT 98.500 120.800 98.900 123.100 ;
        RECT 100.600 120.800 101.000 125.100 ;
        RECT 107.800 120.800 108.200 124.100 ;
        RECT 109.400 120.800 109.800 125.100 ;
        RECT 111.500 120.800 111.900 123.100 ;
        RECT 113.400 120.800 113.900 124.400 ;
        RECT 116.500 121.100 117.000 124.400 ;
        RECT 116.500 120.800 116.900 121.100 ;
        RECT 119.000 120.800 119.400 124.500 ;
        RECT 121.400 120.800 121.800 123.100 ;
        RECT 123.000 120.800 123.400 123.100 ;
        RECT 124.600 120.800 125.000 122.900 ;
        RECT 127.000 120.800 127.500 124.400 ;
        RECT 130.100 121.100 130.600 124.400 ;
        RECT 130.100 120.800 130.500 121.100 ;
        RECT 131.800 120.800 132.200 123.100 ;
        RECT 133.400 120.800 133.800 122.900 ;
        RECT 136.600 120.800 137.000 124.500 ;
        RECT 138.200 120.800 138.600 125.100 ;
        RECT 140.300 120.800 140.700 123.100 ;
        RECT 142.200 120.800 142.700 124.400 ;
        RECT 145.300 121.100 145.800 124.400 ;
        RECT 145.300 120.800 145.700 121.100 ;
        RECT 147.000 120.800 147.400 125.100 ;
        RECT 0.200 120.200 151.800 120.800 ;
        RECT 0.600 117.900 1.000 120.200 ;
        RECT 2.200 117.900 2.600 120.200 ;
        RECT 3.800 116.600 4.300 120.200 ;
        RECT 6.900 119.900 7.300 120.200 ;
        RECT 6.900 116.600 7.400 119.900 ;
        RECT 8.600 115.900 9.000 120.200 ;
        RECT 11.800 116.600 12.300 120.200 ;
        RECT 14.900 119.900 15.300 120.200 ;
        RECT 14.900 116.600 15.400 119.900 ;
        RECT 16.600 117.900 17.000 120.200 ;
        RECT 18.200 115.900 18.600 120.200 ;
        RECT 20.300 117.900 20.700 120.200 ;
        RECT 21.400 117.900 21.800 120.200 ;
        RECT 23.000 117.900 23.400 120.200 ;
        RECT 24.600 116.600 25.100 120.200 ;
        RECT 27.700 119.900 28.100 120.200 ;
        RECT 27.700 116.600 28.200 119.900 ;
        RECT 30.200 116.000 30.600 120.200 ;
        RECT 33.000 117.900 33.400 120.200 ;
        RECT 34.600 117.900 35.000 120.200 ;
        RECT 37.400 115.900 37.800 120.200 ;
        RECT 40.600 115.900 41.000 120.200 ;
        RECT 41.400 117.900 41.800 120.200 ;
        RECT 43.000 117.900 43.400 120.200 ;
        RECT 44.600 115.900 45.000 120.200 ;
        RECT 47.000 115.900 47.400 120.200 ;
        RECT 51.000 115.900 51.400 120.200 ;
        RECT 53.100 117.900 53.500 120.200 ;
        RECT 54.200 117.900 54.600 120.200 ;
        RECT 55.800 117.900 56.200 120.200 ;
        RECT 56.600 115.900 57.000 120.200 ;
        RECT 59.000 115.900 59.400 120.200 ;
        RECT 62.200 117.900 62.600 120.200 ;
        RECT 63.800 116.000 64.200 120.200 ;
        RECT 66.600 117.900 67.000 120.200 ;
        RECT 68.200 117.900 68.600 120.200 ;
        RECT 71.000 115.900 71.400 120.200 ;
        RECT 73.500 119.900 73.900 120.200 ;
        RECT 73.400 116.600 73.900 119.900 ;
        RECT 76.500 116.600 77.000 120.200 ;
        RECT 83.000 116.900 83.400 120.200 ;
        RECT 84.600 115.900 85.000 120.200 ;
        RECT 86.700 117.900 87.100 120.200 ;
        RECT 88.600 117.900 89.000 120.200 ;
        RECT 89.400 117.900 89.800 120.200 ;
        RECT 91.000 118.100 91.400 120.200 ;
        RECT 92.600 117.900 93.000 120.200 ;
        RECT 95.000 118.100 95.400 120.200 ;
        RECT 96.600 117.900 97.000 120.200 ;
        RECT 99.000 116.500 99.400 120.200 ;
        RECT 103.000 116.500 103.400 120.200 ;
        RECT 106.200 116.900 106.600 120.200 ;
        RECT 111.800 115.900 112.200 120.200 ;
        RECT 113.900 117.900 114.300 120.200 ;
        RECT 115.900 119.900 116.300 120.200 ;
        RECT 115.800 116.600 116.300 119.900 ;
        RECT 118.900 116.600 119.400 120.200 ;
        RECT 120.600 117.900 121.000 120.200 ;
        RECT 122.200 118.100 122.600 120.200 ;
        RECT 124.600 118.100 125.000 120.200 ;
        RECT 126.200 117.900 126.600 120.200 ;
        RECT 127.800 116.500 128.200 120.200 ;
        RECT 131.000 116.600 131.500 120.200 ;
        RECT 134.100 119.900 134.500 120.200 ;
        RECT 134.100 116.600 134.600 119.900 ;
        RECT 136.600 118.100 137.000 120.200 ;
        RECT 138.200 117.900 138.600 120.200 ;
        RECT 139.800 116.500 140.200 120.200 ;
        RECT 143.000 118.100 143.400 120.200 ;
        RECT 144.600 117.900 145.000 120.200 ;
        RECT 146.200 117.900 146.600 120.200 ;
        RECT 148.600 116.500 149.000 120.200 ;
        RECT 0.600 100.800 1.000 105.100 ;
        RECT 3.000 100.800 3.400 103.100 ;
        RECT 4.600 100.800 5.000 103.100 ;
        RECT 7.800 100.800 8.200 105.100 ;
        RECT 8.600 100.800 9.000 103.100 ;
        RECT 10.200 100.800 10.600 103.100 ;
        RECT 11.800 100.800 12.200 105.000 ;
        RECT 14.600 100.800 15.000 103.100 ;
        RECT 16.200 100.800 16.600 103.100 ;
        RECT 19.000 100.800 19.400 105.100 ;
        RECT 21.400 100.800 21.800 105.000 ;
        RECT 24.200 100.800 24.600 103.100 ;
        RECT 25.800 100.800 26.200 103.100 ;
        RECT 28.600 100.800 29.000 105.100 ;
        RECT 31.000 101.100 31.500 104.400 ;
        RECT 31.100 100.800 31.500 101.100 ;
        RECT 34.100 100.800 34.600 104.400 ;
        RECT 35.800 100.800 36.200 103.100 ;
        RECT 37.400 100.800 37.800 103.100 ;
        RECT 39.000 100.800 39.500 104.400 ;
        RECT 42.100 101.100 42.600 104.400 ;
        RECT 42.100 100.800 42.500 101.100 ;
        RECT 43.800 100.800 44.200 103.100 ;
        RECT 45.700 100.800 46.100 103.100 ;
        RECT 47.800 100.800 48.200 105.100 ;
        RECT 51.000 100.800 51.500 104.400 ;
        RECT 54.100 101.100 54.600 104.400 ;
        RECT 54.100 100.800 54.500 101.100 ;
        RECT 56.600 100.800 57.000 105.000 ;
        RECT 59.400 100.800 59.800 103.100 ;
        RECT 61.000 100.800 61.400 103.100 ;
        RECT 63.800 100.800 64.200 105.100 ;
        RECT 66.200 100.800 66.600 105.000 ;
        RECT 69.000 100.800 69.400 103.100 ;
        RECT 70.600 100.800 71.000 103.100 ;
        RECT 73.400 100.800 73.800 105.100 ;
        RECT 75.800 101.100 76.300 104.400 ;
        RECT 75.900 100.800 76.300 101.100 ;
        RECT 78.900 100.800 79.400 104.400 ;
        RECT 80.600 100.800 81.000 103.100 ;
        RECT 82.200 100.800 82.600 103.100 ;
        RECT 83.800 100.800 84.200 104.500 ;
        RECT 87.000 100.800 87.400 102.900 ;
        RECT 88.600 100.800 89.000 103.100 ;
        RECT 90.200 100.800 90.600 102.900 ;
        RECT 91.800 100.800 92.200 103.100 ;
        RECT 94.200 100.800 94.600 104.500 ;
        RECT 96.600 100.800 97.000 104.500 ;
        RECT 99.000 100.800 99.400 103.100 ;
        RECT 100.600 100.800 101.000 103.100 ;
        RECT 103.800 100.800 104.200 102.900 ;
        RECT 105.400 100.800 105.800 103.100 ;
        RECT 107.000 100.800 107.400 102.900 ;
        RECT 108.600 100.800 109.000 103.100 ;
        RECT 109.400 100.800 109.800 103.100 ;
        RECT 111.300 100.800 111.700 103.100 ;
        RECT 113.400 100.800 113.800 105.100 ;
        RECT 114.200 100.800 114.600 105.100 ;
        RECT 116.300 100.800 116.700 103.100 ;
        RECT 118.200 100.800 118.600 102.900 ;
        RECT 119.800 100.800 120.200 103.100 ;
        RECT 121.400 100.800 121.800 104.500 ;
        RECT 123.800 100.800 124.200 105.100 ;
        RECT 125.900 100.800 126.300 103.100 ;
        RECT 127.800 100.800 128.200 102.900 ;
        RECT 129.400 100.800 129.800 103.100 ;
        RECT 131.000 100.800 131.400 104.500 ;
        RECT 135.000 100.800 135.400 104.500 ;
        RECT 137.400 100.800 137.900 104.400 ;
        RECT 140.500 101.100 141.000 104.400 ;
        RECT 140.500 100.800 140.900 101.100 ;
        RECT 142.200 100.800 142.600 105.100 ;
        RECT 144.300 100.800 144.700 103.100 ;
        RECT 146.200 100.800 146.600 102.900 ;
        RECT 147.800 100.800 148.200 103.100 ;
        RECT 149.400 100.800 149.800 104.500 ;
        RECT 0.200 100.200 151.800 100.800 ;
        RECT 0.600 97.900 1.000 100.200 ;
        RECT 2.200 97.900 2.600 100.200 ;
        RECT 3.800 97.900 4.200 100.200 ;
        RECT 4.600 95.900 5.000 100.200 ;
        RECT 7.000 97.900 7.400 100.200 ;
        RECT 8.600 97.900 9.000 100.200 ;
        RECT 10.200 96.100 10.600 100.200 ;
        RECT 12.600 96.600 13.100 100.200 ;
        RECT 15.700 99.900 16.100 100.200 ;
        RECT 15.700 96.600 16.200 99.900 ;
        RECT 18.200 96.000 18.600 100.200 ;
        RECT 21.000 97.900 21.400 100.200 ;
        RECT 22.600 97.900 23.000 100.200 ;
        RECT 25.400 95.900 25.800 100.200 ;
        RECT 27.800 96.000 28.200 100.200 ;
        RECT 30.600 97.900 31.000 100.200 ;
        RECT 32.200 97.900 32.600 100.200 ;
        RECT 35.000 95.900 35.400 100.200 ;
        RECT 36.600 95.900 37.000 100.200 ;
        RECT 39.000 97.900 39.400 100.200 ;
        RECT 40.600 97.900 41.000 100.200 ;
        RECT 42.200 96.000 42.600 100.200 ;
        RECT 45.000 97.900 45.400 100.200 ;
        RECT 46.600 97.900 47.000 100.200 ;
        RECT 49.400 95.900 49.800 100.200 ;
        RECT 52.600 95.900 53.000 100.200 ;
        RECT 55.800 97.900 56.200 100.200 ;
        RECT 58.200 96.500 58.600 100.200 ;
        RECT 59.800 97.900 60.200 100.200 ;
        RECT 61.400 98.100 61.800 100.200 ;
        RECT 63.000 95.900 63.400 100.200 ;
        RECT 65.400 95.900 65.800 100.200 ;
        RECT 68.600 95.900 69.000 100.200 ;
        RECT 69.400 95.900 69.800 100.200 ;
        RECT 71.500 97.900 71.900 100.200 ;
        RECT 72.600 95.900 73.000 100.200 ;
        RECT 74.700 97.900 75.100 100.200 ;
        RECT 76.600 97.900 77.000 100.200 ;
        RECT 77.700 97.900 78.100 100.200 ;
        RECT 79.800 95.900 80.200 100.200 ;
        RECT 80.600 95.900 81.000 100.200 ;
        RECT 82.700 97.900 83.100 100.200 ;
        RECT 83.800 97.900 84.200 100.200 ;
        RECT 85.400 97.900 85.800 100.200 ;
        RECT 86.200 97.900 86.600 100.200 ;
        RECT 87.800 97.900 88.200 100.200 ;
        RECT 88.600 97.900 89.000 100.200 ;
        RECT 90.200 97.900 90.600 100.200 ;
        RECT 91.000 97.900 91.400 100.200 ;
        RECT 92.600 98.100 93.000 100.200 ;
        RECT 94.200 97.900 94.600 100.200 ;
        RECT 95.800 97.900 96.200 100.200 ;
        RECT 96.600 97.900 97.000 100.200 ;
        RECT 98.200 97.900 98.600 100.200 ;
        RECT 100.600 95.900 101.000 100.200 ;
        RECT 103.800 95.900 104.200 100.200 ;
        RECT 105.400 96.500 105.800 100.200 ;
        RECT 108.600 97.900 109.000 100.200 ;
        RECT 110.200 97.900 110.600 100.200 ;
        RECT 111.000 97.900 111.400 100.200 ;
        RECT 112.600 98.100 113.000 100.200 ;
        RECT 115.000 96.500 115.400 100.200 ;
        RECT 119.000 95.900 119.400 100.200 ;
        RECT 119.800 95.900 120.200 100.200 ;
        RECT 121.900 97.900 122.300 100.200 ;
        RECT 123.000 97.900 123.400 100.200 ;
        RECT 124.600 98.100 125.000 100.200 ;
        RECT 127.000 98.100 127.400 100.200 ;
        RECT 128.600 97.900 129.000 100.200 ;
        RECT 130.200 98.100 130.600 100.200 ;
        RECT 131.800 97.900 132.200 100.200 ;
        RECT 133.400 98.100 133.800 100.200 ;
        RECT 135.000 97.900 135.400 100.200 ;
        RECT 135.800 97.900 136.200 100.200 ;
        RECT 137.400 98.100 137.800 100.200 ;
        RECT 139.000 97.900 139.400 100.200 ;
        RECT 140.600 98.100 141.000 100.200 ;
        RECT 143.000 96.500 143.400 100.200 ;
        RECT 145.400 97.900 145.800 100.200 ;
        RECT 147.000 97.900 147.400 100.200 ;
        RECT 148.600 98.100 149.000 100.200 ;
        RECT 150.200 97.900 150.600 100.200 ;
        RECT 0.600 80.800 1.000 83.100 ;
        RECT 2.200 80.800 2.600 83.100 ;
        RECT 3.800 80.800 4.200 83.100 ;
        RECT 5.900 80.800 6.300 85.100 ;
        RECT 7.800 80.800 8.200 83.100 ;
        RECT 9.400 80.800 9.800 84.900 ;
        RECT 11.300 80.800 11.700 83.100 ;
        RECT 13.400 80.800 13.800 85.100 ;
        RECT 14.200 80.800 14.600 83.100 ;
        RECT 17.400 80.800 17.800 84.500 ;
        RECT 19.000 80.800 19.400 85.100 ;
        RECT 21.400 80.800 21.800 85.100 ;
        RECT 23.800 80.800 24.300 84.400 ;
        RECT 26.900 81.100 27.400 84.400 ;
        RECT 26.900 80.800 27.300 81.100 ;
        RECT 29.400 80.800 29.800 85.000 ;
        RECT 32.200 80.800 32.600 83.100 ;
        RECT 33.800 80.800 34.200 83.100 ;
        RECT 36.600 80.800 37.000 85.100 ;
        RECT 39.000 80.800 39.400 85.000 ;
        RECT 41.800 80.800 42.200 83.100 ;
        RECT 43.400 80.800 43.800 83.100 ;
        RECT 46.200 80.800 46.600 85.100 ;
        RECT 50.200 80.800 50.600 85.000 ;
        RECT 53.000 80.800 53.400 83.100 ;
        RECT 54.600 80.800 55.000 83.100 ;
        RECT 57.400 80.800 57.800 85.100 ;
        RECT 59.000 80.800 59.400 83.100 ;
        RECT 60.600 80.800 61.000 83.100 ;
        RECT 62.200 80.800 62.600 84.900 ;
        RECT 63.800 80.800 64.200 83.100 ;
        RECT 65.400 80.800 65.800 83.100 ;
        RECT 66.200 80.800 66.600 83.100 ;
        RECT 67.800 80.800 68.200 83.100 ;
        RECT 68.600 80.800 69.000 83.100 ;
        RECT 70.200 80.800 70.600 83.100 ;
        RECT 73.400 80.800 73.800 84.500 ;
        RECT 75.000 80.800 75.400 83.100 ;
        RECT 76.600 80.800 77.000 83.100 ;
        RECT 77.400 80.800 77.800 83.100 ;
        RECT 79.000 80.800 79.400 83.100 ;
        RECT 81.400 80.800 81.800 84.500 ;
        RECT 83.800 80.800 84.200 83.100 ;
        RECT 85.400 80.800 85.800 84.500 ;
        RECT 87.800 80.800 88.200 83.100 ;
        RECT 89.400 80.800 89.800 83.100 ;
        RECT 90.200 80.800 90.600 83.100 ;
        RECT 91.800 80.800 92.200 85.100 ;
        RECT 93.900 80.800 94.300 83.100 ;
        RECT 97.400 80.800 97.800 84.500 ;
        RECT 99.000 80.800 99.400 83.100 ;
        RECT 100.600 80.800 101.000 83.100 ;
        RECT 103.000 80.800 103.400 83.100 ;
        RECT 104.600 80.800 105.000 83.100 ;
        RECT 105.400 80.800 105.800 83.100 ;
        RECT 107.000 80.800 107.400 82.900 ;
        RECT 109.400 80.800 109.800 84.500 ;
        RECT 111.800 80.800 112.200 83.100 ;
        RECT 113.400 80.800 113.800 82.900 ;
        RECT 115.800 80.800 116.200 84.500 ;
        RECT 118.200 80.800 118.600 85.100 ;
        RECT 121.400 80.800 121.800 85.100 ;
        RECT 122.200 80.800 122.600 85.100 ;
        RECT 124.900 80.800 125.300 83.100 ;
        RECT 127.000 80.800 127.400 85.100 ;
        RECT 127.800 80.800 128.200 85.100 ;
        RECT 129.900 80.800 130.300 83.100 ;
        RECT 132.600 80.800 133.000 84.500 ;
        RECT 135.000 80.800 135.400 82.900 ;
        RECT 136.600 80.800 137.000 83.100 ;
        RECT 138.200 80.800 138.600 82.900 ;
        RECT 139.800 80.800 140.200 83.100 ;
        RECT 141.400 80.800 141.800 84.500 ;
        RECT 143.800 80.800 144.200 83.100 ;
        RECT 145.400 80.800 145.800 82.900 ;
        RECT 147.000 80.800 147.400 83.100 ;
        RECT 148.600 80.800 149.000 82.900 ;
        RECT 0.200 80.200 151.800 80.800 ;
        RECT 0.600 77.900 1.000 80.200 ;
        RECT 2.200 77.900 2.600 80.200 ;
        RECT 3.800 75.900 4.200 80.200 ;
        RECT 7.100 79.900 7.500 80.200 ;
        RECT 7.000 76.600 7.500 79.900 ;
        RECT 10.100 76.600 10.600 80.200 ;
        RECT 11.800 77.900 12.200 80.200 ;
        RECT 13.400 75.900 13.800 80.200 ;
        RECT 15.500 77.900 15.900 80.200 ;
        RECT 18.200 76.500 18.600 80.200 ;
        RECT 20.600 76.000 21.000 80.200 ;
        RECT 23.400 77.900 23.800 80.200 ;
        RECT 25.000 77.900 25.400 80.200 ;
        RECT 27.800 75.900 28.200 80.200 ;
        RECT 30.200 76.000 30.600 80.200 ;
        RECT 33.000 77.900 33.400 80.200 ;
        RECT 34.600 77.900 35.000 80.200 ;
        RECT 37.400 75.900 37.800 80.200 ;
        RECT 39.800 76.000 40.200 80.200 ;
        RECT 42.600 77.900 43.000 80.200 ;
        RECT 44.200 77.900 44.600 80.200 ;
        RECT 47.000 75.900 47.400 80.200 ;
        RECT 51.000 76.000 51.400 80.200 ;
        RECT 53.800 77.900 54.200 80.200 ;
        RECT 55.400 77.900 55.800 80.200 ;
        RECT 58.200 75.900 58.600 80.200 ;
        RECT 59.800 77.900 60.200 80.200 ;
        RECT 61.400 77.900 61.800 80.200 ;
        RECT 63.000 78.100 63.400 80.200 ;
        RECT 64.600 77.900 65.000 80.200 ;
        RECT 67.000 76.500 67.400 80.200 ;
        RECT 68.600 77.900 69.000 80.200 ;
        RECT 70.200 77.900 70.600 80.200 ;
        RECT 72.600 76.500 73.000 80.200 ;
        RECT 75.000 76.500 75.400 80.200 ;
        RECT 76.600 75.900 77.000 80.200 ;
        RECT 78.200 76.500 78.600 80.200 ;
        RECT 79.800 75.900 80.200 80.200 ;
        RECT 81.400 76.500 81.800 80.200 ;
        RECT 83.000 75.900 83.400 80.200 ;
        RECT 83.800 77.900 84.200 80.200 ;
        RECT 85.400 77.900 85.800 80.200 ;
        RECT 87.000 76.500 87.400 80.200 ;
        RECT 90.200 77.900 90.600 80.200 ;
        RECT 91.800 77.900 92.200 80.200 ;
        RECT 95.000 76.500 95.400 80.200 ;
        RECT 97.400 76.500 97.800 80.200 ;
        RECT 102.200 76.500 102.600 80.200 ;
        RECT 104.600 77.900 105.000 80.200 ;
        RECT 106.200 77.900 106.600 80.200 ;
        RECT 107.000 75.900 107.400 80.200 ;
        RECT 109.400 77.900 109.800 80.200 ;
        RECT 111.000 77.900 111.400 80.200 ;
        RECT 112.600 78.100 113.000 80.200 ;
        RECT 114.200 77.900 114.600 80.200 ;
        RECT 115.800 78.100 116.200 80.200 ;
        RECT 117.400 77.900 117.800 80.200 ;
        RECT 119.000 75.900 119.400 80.200 ;
        RECT 119.800 77.900 120.200 80.200 ;
        RECT 121.400 78.100 121.800 80.200 ;
        RECT 123.800 76.500 124.200 80.200 ;
        RECT 126.200 77.900 126.600 80.200 ;
        RECT 127.800 78.100 128.200 80.200 ;
        RECT 129.400 75.900 129.800 80.200 ;
        RECT 131.500 77.900 131.900 80.200 ;
        RECT 133.500 79.900 133.900 80.200 ;
        RECT 133.400 76.600 133.900 79.900 ;
        RECT 136.500 76.600 137.000 80.200 ;
        RECT 138.200 77.900 138.600 80.200 ;
        RECT 139.800 78.100 140.200 80.200 ;
        RECT 141.400 77.900 141.800 80.200 ;
        RECT 143.000 78.100 143.400 80.200 ;
        RECT 145.400 78.100 145.800 80.200 ;
        RECT 147.000 77.900 147.400 80.200 ;
        RECT 148.600 76.500 149.000 80.200 ;
        RECT 0.600 60.800 1.000 65.100 ;
        RECT 3.800 60.800 4.300 64.400 ;
        RECT 6.900 61.100 7.400 64.400 ;
        RECT 6.900 60.800 7.300 61.100 ;
        RECT 8.600 60.800 9.000 63.100 ;
        RECT 11.000 60.800 11.400 64.500 ;
        RECT 15.000 60.800 15.400 65.100 ;
        RECT 15.800 60.800 16.200 63.100 ;
        RECT 17.400 60.800 17.800 63.100 ;
        RECT 19.000 60.800 19.500 64.400 ;
        RECT 22.100 61.100 22.600 64.400 ;
        RECT 22.100 60.800 22.500 61.100 ;
        RECT 24.600 60.800 25.100 64.400 ;
        RECT 27.700 61.100 28.200 64.400 ;
        RECT 27.700 60.800 28.100 61.100 ;
        RECT 30.200 60.800 30.700 64.400 ;
        RECT 33.300 61.100 33.800 64.400 ;
        RECT 33.300 60.800 33.700 61.100 ;
        RECT 35.000 60.800 35.400 65.100 ;
        RECT 38.200 60.800 38.600 65.000 ;
        RECT 41.000 60.800 41.400 63.100 ;
        RECT 42.600 60.800 43.000 63.100 ;
        RECT 45.400 60.800 45.800 65.100 ;
        RECT 49.400 60.800 49.800 65.000 ;
        RECT 52.200 60.800 52.600 63.100 ;
        RECT 53.800 60.800 54.200 63.100 ;
        RECT 56.600 60.800 57.000 65.100 ;
        RECT 58.200 60.800 58.600 63.100 ;
        RECT 59.800 60.800 60.200 63.100 ;
        RECT 60.600 60.800 61.000 63.100 ;
        RECT 62.200 60.800 62.600 63.100 ;
        RECT 63.800 60.800 64.200 62.900 ;
        RECT 65.400 60.800 65.800 63.100 ;
        RECT 67.000 60.800 67.400 62.900 ;
        RECT 68.600 60.800 69.000 63.100 ;
        RECT 69.400 60.800 69.800 63.100 ;
        RECT 71.300 60.800 71.700 63.100 ;
        RECT 73.400 60.800 73.800 65.100 ;
        RECT 74.200 60.800 74.600 65.100 ;
        RECT 76.300 60.800 76.700 63.100 ;
        RECT 77.400 60.800 77.800 63.100 ;
        RECT 79.000 60.800 79.400 63.100 ;
        RECT 79.800 60.800 80.200 63.100 ;
        RECT 81.400 60.800 81.800 63.100 ;
        RECT 82.200 60.800 82.600 65.100 ;
        RECT 83.800 60.800 84.200 64.500 ;
        RECT 86.200 60.800 86.600 64.500 ;
        RECT 87.800 60.800 88.200 65.100 ;
        RECT 88.600 60.800 89.000 63.100 ;
        RECT 90.200 60.800 90.600 63.100 ;
        RECT 91.000 60.800 91.400 65.100 ;
        RECT 94.200 60.800 94.600 65.100 ;
        RECT 95.300 60.800 95.700 63.100 ;
        RECT 97.400 60.800 97.800 65.100 ;
        RECT 98.200 60.800 98.600 65.100 ;
        RECT 100.300 60.800 100.700 63.100 ;
        RECT 103.000 60.800 103.400 65.100 ;
        RECT 104.900 60.800 105.300 63.100 ;
        RECT 107.000 60.800 107.400 65.100 ;
        RECT 107.800 60.800 108.200 65.100 ;
        RECT 109.900 60.800 110.300 63.100 ;
        RECT 111.800 60.800 112.200 64.500 ;
        RECT 114.200 60.800 114.600 63.100 ;
        RECT 115.800 60.800 116.200 62.900 ;
        RECT 118.200 60.800 118.600 62.900 ;
        RECT 119.800 60.800 120.200 63.100 ;
        RECT 120.600 60.800 121.000 63.100 ;
        RECT 122.200 60.800 122.600 62.900 ;
        RECT 124.600 60.800 125.000 64.500 ;
        RECT 127.000 60.800 127.400 63.100 ;
        RECT 128.600 60.800 129.000 62.900 ;
        RECT 130.200 60.800 130.600 63.100 ;
        RECT 131.800 60.800 132.200 62.900 ;
        RECT 133.400 60.800 133.800 63.100 ;
        RECT 135.000 60.800 135.400 62.900 ;
        RECT 137.400 60.800 137.800 64.500 ;
        RECT 140.600 60.800 141.000 62.900 ;
        RECT 142.200 60.800 142.600 63.100 ;
        RECT 143.800 60.800 144.200 62.900 ;
        RECT 145.400 60.800 145.800 63.100 ;
        RECT 147.000 60.800 147.500 64.400 ;
        RECT 150.100 61.100 150.600 64.400 ;
        RECT 150.100 60.800 150.500 61.100 ;
        RECT 0.200 60.200 151.800 60.800 ;
        RECT 1.500 59.900 1.900 60.200 ;
        RECT 1.400 56.600 1.900 59.900 ;
        RECT 4.500 56.600 5.000 60.200 ;
        RECT 7.000 56.000 7.400 60.200 ;
        RECT 9.800 57.900 10.200 60.200 ;
        RECT 11.400 57.900 11.800 60.200 ;
        RECT 14.200 55.900 14.600 60.200 ;
        RECT 16.700 59.900 17.100 60.200 ;
        RECT 16.600 56.600 17.100 59.900 ;
        RECT 19.700 56.600 20.200 60.200 ;
        RECT 21.400 57.900 21.800 60.200 ;
        RECT 23.000 57.900 23.400 60.200 ;
        RECT 23.800 57.900 24.200 60.200 ;
        RECT 25.400 55.900 25.800 60.200 ;
        RECT 27.800 55.900 28.200 60.200 ;
        RECT 30.200 57.900 30.600 60.200 ;
        RECT 31.800 55.900 32.200 60.200 ;
        RECT 33.400 55.900 33.800 60.200 ;
        RECT 35.000 55.900 35.400 60.200 ;
        RECT 36.600 55.900 37.000 60.200 ;
        RECT 38.200 55.900 38.600 60.200 ;
        RECT 39.800 56.000 40.200 60.200 ;
        RECT 42.600 57.900 43.000 60.200 ;
        RECT 44.200 57.900 44.600 60.200 ;
        RECT 47.000 55.900 47.400 60.200 ;
        RECT 51.000 56.500 51.400 60.200 ;
        RECT 54.200 58.100 54.600 60.200 ;
        RECT 55.800 57.900 56.200 60.200 ;
        RECT 56.600 57.900 57.000 60.200 ;
        RECT 58.200 57.900 58.600 60.200 ;
        RECT 59.000 57.900 59.400 60.200 ;
        RECT 60.600 57.900 61.000 60.200 ;
        RECT 61.400 57.900 61.800 60.200 ;
        RECT 63.000 57.900 63.400 60.200 ;
        RECT 63.800 57.900 64.200 60.200 ;
        RECT 65.400 57.900 65.800 60.200 ;
        RECT 67.000 56.500 67.400 60.200 ;
        RECT 68.600 55.900 69.000 60.200 ;
        RECT 69.400 55.900 69.800 60.200 ;
        RECT 71.500 57.900 71.900 60.200 ;
        RECT 72.600 57.900 73.000 60.200 ;
        RECT 74.200 57.900 74.600 60.200 ;
        RECT 75.000 57.900 75.400 60.200 ;
        RECT 76.600 57.900 77.000 60.200 ;
        RECT 77.400 57.900 77.800 60.200 ;
        RECT 79.000 57.900 79.400 60.200 ;
        RECT 79.800 57.900 80.200 60.200 ;
        RECT 81.400 57.900 81.800 60.200 ;
        RECT 82.200 55.900 82.600 60.200 ;
        RECT 84.600 55.900 85.000 60.200 ;
        RECT 87.800 55.900 88.200 60.200 ;
        RECT 90.200 56.500 90.600 60.200 ;
        RECT 91.800 57.900 92.200 60.200 ;
        RECT 93.400 58.100 93.800 60.200 ;
        RECT 95.800 58.100 96.200 60.200 ;
        RECT 97.400 57.900 97.800 60.200 ;
        RECT 99.000 56.500 99.400 60.200 ;
        RECT 103.000 55.900 103.400 60.200 ;
        RECT 105.100 57.900 105.500 60.200 ;
        RECT 107.000 58.100 107.400 60.200 ;
        RECT 108.600 57.900 109.000 60.200 ;
        RECT 110.200 56.500 110.600 60.200 ;
        RECT 112.600 57.900 113.000 60.200 ;
        RECT 114.200 58.100 114.600 60.200 ;
        RECT 116.600 58.100 117.000 60.200 ;
        RECT 118.200 57.900 118.600 60.200 ;
        RECT 119.800 56.500 120.200 60.200 ;
        RECT 123.000 58.100 123.400 60.200 ;
        RECT 124.600 57.900 125.000 60.200 ;
        RECT 127.000 56.500 127.400 60.200 ;
        RECT 128.600 55.900 129.000 60.200 ;
        RECT 130.700 57.900 131.100 60.200 ;
        RECT 132.600 58.100 133.000 60.200 ;
        RECT 134.200 57.900 134.600 60.200 ;
        RECT 135.000 57.900 135.400 60.200 ;
        RECT 136.600 58.100 137.000 60.200 ;
        RECT 138.200 57.900 138.600 60.200 ;
        RECT 139.800 57.900 140.200 60.200 ;
        RECT 141.400 55.900 141.800 60.200 ;
        RECT 143.000 56.600 143.500 60.200 ;
        RECT 146.100 59.900 146.500 60.200 ;
        RECT 146.100 56.600 146.600 59.900 ;
        RECT 147.800 55.900 148.200 60.200 ;
        RECT 149.900 57.900 150.300 60.200 ;
        RECT 0.600 40.800 1.000 43.100 ;
        RECT 2.200 40.800 2.600 43.100 ;
        RECT 3.800 40.800 4.300 44.400 ;
        RECT 6.900 41.100 7.400 44.400 ;
        RECT 6.900 40.800 7.300 41.100 ;
        RECT 8.900 40.800 9.300 43.100 ;
        RECT 11.000 40.800 11.400 45.100 ;
        RECT 12.600 40.800 13.100 44.400 ;
        RECT 15.700 41.100 16.200 44.400 ;
        RECT 15.700 40.800 16.100 41.100 ;
        RECT 18.200 40.800 18.600 45.000 ;
        RECT 21.000 40.800 21.400 43.100 ;
        RECT 22.600 40.800 23.000 43.100 ;
        RECT 25.400 40.800 25.800 45.100 ;
        RECT 27.000 40.800 27.400 45.100 ;
        RECT 28.600 40.800 29.000 45.100 ;
        RECT 30.200 40.800 30.600 45.100 ;
        RECT 31.800 40.800 32.200 45.100 ;
        RECT 33.400 40.800 33.800 45.100 ;
        RECT 35.800 40.800 36.200 45.100 ;
        RECT 36.600 40.800 37.000 43.100 ;
        RECT 38.200 40.800 38.600 44.900 ;
        RECT 39.800 40.800 40.200 45.100 ;
        RECT 41.900 40.800 42.300 43.100 ;
        RECT 43.800 40.800 44.200 43.100 ;
        RECT 44.600 40.800 45.000 45.100 ;
        RECT 48.600 40.800 49.000 44.500 ;
        RECT 52.600 40.800 53.100 44.400 ;
        RECT 55.700 41.100 56.200 44.400 ;
        RECT 55.700 40.800 56.100 41.100 ;
        RECT 58.200 40.800 58.600 45.000 ;
        RECT 61.000 40.800 61.400 43.100 ;
        RECT 62.600 40.800 63.000 43.100 ;
        RECT 65.400 40.800 65.800 45.100 ;
        RECT 67.000 40.800 67.400 45.100 ;
        RECT 68.600 40.800 69.000 45.100 ;
        RECT 70.200 40.800 70.600 45.100 ;
        RECT 71.800 40.800 72.200 45.100 ;
        RECT 73.400 40.800 73.800 45.100 ;
        RECT 74.200 40.800 74.600 45.100 ;
        RECT 76.900 40.800 77.300 43.100 ;
        RECT 79.000 40.800 79.400 45.100 ;
        RECT 80.600 40.800 81.000 43.100 ;
        RECT 81.700 40.800 82.100 43.100 ;
        RECT 83.800 40.800 84.200 45.100 ;
        RECT 84.600 40.800 85.000 45.100 ;
        RECT 86.200 40.800 86.600 45.100 ;
        RECT 88.600 40.800 89.000 45.100 ;
        RECT 91.800 40.800 92.200 44.500 ;
        RECT 93.400 40.800 93.800 45.100 ;
        RECT 94.200 40.800 94.600 45.100 ;
        RECT 96.100 40.800 96.500 43.100 ;
        RECT 98.200 40.800 98.600 45.100 ;
        RECT 100.600 40.800 101.000 45.100 ;
        RECT 104.600 40.800 105.000 44.500 ;
        RECT 107.000 40.800 107.400 43.100 ;
        RECT 107.800 40.800 108.200 45.100 ;
        RECT 109.900 40.800 110.300 43.100 ;
        RECT 111.000 40.800 111.400 45.100 ;
        RECT 113.100 40.800 113.500 43.100 ;
        RECT 114.200 40.800 114.600 43.100 ;
        RECT 117.400 40.800 117.800 44.500 ;
        RECT 119.000 40.800 119.400 43.100 ;
        RECT 120.600 40.800 121.000 42.900 ;
        RECT 122.200 40.800 122.600 45.100 ;
        RECT 124.600 40.800 125.000 44.500 ;
        RECT 127.000 40.800 127.400 45.100 ;
        RECT 129.100 40.800 129.500 43.100 ;
        RECT 131.000 40.800 131.400 42.900 ;
        RECT 132.600 40.800 133.000 43.100 ;
        RECT 135.000 40.800 135.400 44.500 ;
        RECT 137.900 40.800 138.300 45.100 ;
        RECT 139.800 40.800 140.200 43.100 ;
        RECT 141.400 40.800 141.800 43.100 ;
        RECT 142.200 40.800 142.600 43.100 ;
        RECT 143.800 40.800 144.200 42.900 ;
        RECT 145.400 40.800 145.800 45.100 ;
        RECT 147.800 40.800 148.200 43.100 ;
        RECT 149.400 40.800 149.800 44.900 ;
        RECT 0.200 40.200 151.800 40.800 ;
        RECT 1.500 39.900 1.900 40.200 ;
        RECT 1.400 36.600 1.900 39.900 ;
        RECT 4.500 36.600 5.000 40.200 ;
        RECT 6.200 37.900 6.600 40.200 ;
        RECT 7.800 37.900 8.200 40.200 ;
        RECT 9.400 37.900 9.800 40.200 ;
        RECT 10.500 37.900 10.900 40.200 ;
        RECT 12.600 35.900 13.000 40.200 ;
        RECT 14.200 36.600 14.700 40.200 ;
        RECT 17.300 39.900 17.700 40.200 ;
        RECT 17.300 36.600 17.800 39.900 ;
        RECT 19.800 36.000 20.200 40.200 ;
        RECT 22.600 37.900 23.000 40.200 ;
        RECT 24.200 37.900 24.600 40.200 ;
        RECT 27.000 35.900 27.400 40.200 ;
        RECT 29.400 36.000 29.800 40.200 ;
        RECT 32.200 37.900 32.600 40.200 ;
        RECT 33.800 37.900 34.200 40.200 ;
        RECT 36.600 35.900 37.000 40.200 ;
        RECT 39.000 37.900 39.400 40.200 ;
        RECT 40.600 36.600 41.100 40.200 ;
        RECT 43.700 39.900 44.100 40.200 ;
        RECT 43.700 36.600 44.200 39.900 ;
        RECT 45.400 37.900 45.800 40.200 ;
        RECT 47.000 37.900 47.400 40.200 ;
        RECT 50.300 39.900 50.700 40.200 ;
        RECT 50.200 36.600 50.700 39.900 ;
        RECT 53.300 36.600 53.800 40.200 ;
        RECT 55.800 36.000 56.200 40.200 ;
        RECT 58.600 37.900 59.000 40.200 ;
        RECT 60.200 37.900 60.600 40.200 ;
        RECT 63.000 35.900 63.400 40.200 ;
        RECT 65.400 36.000 65.800 40.200 ;
        RECT 68.200 37.900 68.600 40.200 ;
        RECT 69.800 37.900 70.200 40.200 ;
        RECT 72.600 35.900 73.000 40.200 ;
        RECT 74.200 35.900 74.600 40.200 ;
        RECT 75.800 35.900 76.200 40.200 ;
        RECT 78.200 35.900 78.600 40.200 ;
        RECT 79.000 37.900 79.400 40.200 ;
        RECT 80.600 35.900 81.000 40.200 ;
        RECT 82.700 37.900 83.100 40.200 ;
        RECT 85.400 35.900 85.800 40.200 ;
        RECT 86.500 37.900 86.900 40.200 ;
        RECT 88.600 35.900 89.000 40.200 ;
        RECT 89.700 37.900 90.100 40.200 ;
        RECT 91.800 35.900 92.200 40.200 ;
        RECT 93.400 37.900 93.800 40.200 ;
        RECT 95.000 36.500 95.400 40.200 ;
        RECT 96.600 35.900 97.000 40.200 ;
        RECT 97.400 35.900 97.800 40.200 ;
        RECT 99.500 37.900 99.900 40.200 ;
        RECT 102.200 37.900 102.600 40.200 ;
        RECT 103.800 37.900 104.200 40.200 ;
        RECT 104.600 37.900 105.000 40.200 ;
        RECT 107.800 36.500 108.200 40.200 ;
        RECT 109.400 37.900 109.800 40.200 ;
        RECT 111.000 38.100 111.400 40.200 ;
        RECT 112.600 35.900 113.000 40.200 ;
        RECT 114.700 37.900 115.100 40.200 ;
        RECT 117.400 36.500 117.800 40.200 ;
        RECT 119.000 37.900 119.400 40.200 ;
        RECT 120.600 37.900 121.000 40.200 ;
        RECT 121.400 35.900 121.800 40.200 ;
        RECT 123.500 37.900 123.900 40.200 ;
        RECT 126.200 36.500 126.600 40.200 ;
        RECT 128.600 38.100 129.000 40.200 ;
        RECT 130.200 37.900 130.600 40.200 ;
        RECT 131.000 37.900 131.400 40.200 ;
        RECT 132.600 38.100 133.000 40.200 ;
        RECT 135.800 36.500 136.200 40.200 ;
        RECT 138.200 38.100 138.600 40.200 ;
        RECT 139.800 37.900 140.200 40.200 ;
        RECT 141.400 36.500 141.800 40.200 ;
        RECT 143.800 37.900 144.200 40.200 ;
        RECT 145.400 38.100 145.800 40.200 ;
        RECT 147.300 37.900 147.700 40.200 ;
        RECT 149.400 35.900 149.800 40.200 ;
        RECT 0.600 20.800 1.000 25.100 ;
        RECT 2.200 20.800 2.600 25.100 ;
        RECT 3.800 20.800 4.200 25.100 ;
        RECT 5.400 20.800 5.800 25.100 ;
        RECT 7.000 20.800 7.400 25.100 ;
        RECT 8.600 20.800 9.100 24.400 ;
        RECT 11.700 21.100 12.200 24.400 ;
        RECT 11.700 20.800 12.100 21.100 ;
        RECT 14.200 20.800 14.600 25.000 ;
        RECT 17.000 20.800 17.400 23.100 ;
        RECT 18.600 20.800 19.000 23.100 ;
        RECT 21.400 20.800 21.800 25.100 ;
        RECT 23.800 20.800 24.200 25.000 ;
        RECT 26.600 20.800 27.000 23.100 ;
        RECT 28.200 20.800 28.600 23.100 ;
        RECT 31.000 20.800 31.400 25.100 ;
        RECT 33.400 20.800 33.800 25.000 ;
        RECT 36.200 20.800 36.600 23.100 ;
        RECT 37.800 20.800 38.200 23.100 ;
        RECT 40.600 20.800 41.000 25.100 ;
        RECT 43.000 20.800 43.400 25.000 ;
        RECT 45.800 20.800 46.200 23.100 ;
        RECT 47.400 20.800 47.800 23.100 ;
        RECT 50.200 20.800 50.600 25.100 ;
        RECT 54.200 20.800 54.600 25.000 ;
        RECT 57.000 20.800 57.400 23.100 ;
        RECT 58.600 20.800 59.000 23.100 ;
        RECT 61.400 20.800 61.800 25.100 ;
        RECT 63.000 20.800 63.400 25.100 ;
        RECT 64.600 20.800 65.000 25.100 ;
        RECT 66.200 20.800 66.600 25.100 ;
        RECT 67.800 20.800 68.200 25.100 ;
        RECT 69.400 20.800 69.800 25.100 ;
        RECT 70.200 20.800 70.600 25.100 ;
        RECT 71.800 20.800 72.200 25.100 ;
        RECT 73.400 20.800 73.800 25.100 ;
        RECT 75.000 20.800 75.400 25.100 ;
        RECT 76.600 20.800 77.000 25.100 ;
        RECT 78.200 21.100 78.700 24.400 ;
        RECT 78.300 20.800 78.700 21.100 ;
        RECT 81.300 20.800 81.800 24.400 ;
        RECT 83.800 20.800 84.200 23.100 ;
        RECT 86.200 20.800 86.600 24.500 ;
        RECT 89.400 20.800 89.800 25.100 ;
        RECT 90.200 20.800 90.600 23.100 ;
        RECT 92.100 20.800 92.500 23.100 ;
        RECT 94.200 20.800 94.600 25.100 ;
        RECT 96.600 20.800 97.000 24.500 ;
        RECT 99.000 20.800 99.400 22.900 ;
        RECT 100.600 20.800 101.000 23.100 ;
        RECT 104.600 20.800 105.000 24.500 ;
        RECT 107.000 20.800 107.400 22.900 ;
        RECT 108.600 20.800 109.000 23.100 ;
        RECT 110.200 20.800 110.600 23.100 ;
        RECT 111.000 20.800 111.400 25.100 ;
        RECT 114.700 20.800 115.100 25.100 ;
        RECT 121.400 20.800 121.800 24.100 ;
        RECT 123.000 20.800 123.400 25.100 ;
        RECT 125.100 20.800 125.500 23.100 ;
        RECT 126.200 20.800 126.600 25.100 ;
        RECT 129.400 20.800 129.800 24.500 ;
        RECT 134.200 20.800 134.600 25.100 ;
        RECT 135.800 20.800 136.200 22.900 ;
        RECT 137.400 20.800 137.800 23.100 ;
        RECT 138.200 20.800 138.600 25.100 ;
        RECT 140.300 20.800 140.700 23.100 ;
        RECT 141.400 20.800 141.800 23.100 ;
        RECT 143.000 20.800 143.400 23.100 ;
        RECT 143.800 20.800 144.200 23.100 ;
        RECT 145.400 20.800 145.800 22.900 ;
        RECT 147.300 20.800 147.700 23.100 ;
        RECT 149.400 20.800 149.800 25.100 ;
        RECT 0.200 20.200 151.800 20.800 ;
        RECT 1.400 16.000 1.800 20.200 ;
        RECT 4.200 17.900 4.600 20.200 ;
        RECT 5.800 17.900 6.200 20.200 ;
        RECT 8.600 15.900 9.000 20.200 ;
        RECT 10.200 17.900 10.600 20.200 ;
        RECT 12.700 19.900 13.100 20.200 ;
        RECT 12.600 16.600 13.100 19.900 ;
        RECT 15.700 16.600 16.200 20.200 ;
        RECT 18.200 16.000 18.600 20.200 ;
        RECT 21.000 17.900 21.400 20.200 ;
        RECT 22.600 17.900 23.000 20.200 ;
        RECT 25.400 15.900 25.800 20.200 ;
        RECT 27.900 19.900 28.300 20.200 ;
        RECT 27.800 16.600 28.300 19.900 ;
        RECT 30.900 16.600 31.400 20.200 ;
        RECT 33.400 16.000 33.800 20.200 ;
        RECT 36.200 17.900 36.600 20.200 ;
        RECT 37.800 17.900 38.200 20.200 ;
        RECT 40.600 15.900 41.000 20.200 ;
        RECT 43.000 16.100 43.400 20.200 ;
        RECT 44.600 17.900 45.000 20.200 ;
        RECT 47.000 15.900 47.400 20.200 ;
        RECT 47.800 15.900 48.200 20.200 ;
        RECT 52.600 16.000 53.000 20.200 ;
        RECT 55.400 17.900 55.800 20.200 ;
        RECT 57.000 17.900 57.400 20.200 ;
        RECT 59.800 15.900 60.200 20.200 ;
        RECT 62.200 16.000 62.600 20.200 ;
        RECT 65.000 17.900 65.400 20.200 ;
        RECT 66.600 17.900 67.000 20.200 ;
        RECT 69.400 15.900 69.800 20.200 ;
        RECT 71.000 17.900 71.400 20.200 ;
        RECT 72.600 17.900 73.000 20.200 ;
        RECT 75.000 15.900 75.400 20.200 ;
        RECT 75.800 17.900 76.200 20.200 ;
        RECT 77.400 15.900 77.800 20.200 ;
        RECT 79.500 17.900 79.900 20.200 ;
        RECT 82.200 15.900 82.600 20.200 ;
        RECT 83.800 16.100 84.200 20.200 ;
        RECT 85.400 17.900 85.800 20.200 ;
        RECT 87.000 16.100 87.400 20.200 ;
        RECT 88.600 17.900 89.000 20.200 ;
        RECT 90.200 17.900 90.600 20.200 ;
        RECT 92.600 16.500 93.000 20.200 ;
        RECT 94.200 17.900 94.600 20.200 ;
        RECT 95.800 18.100 96.200 20.200 ;
        RECT 97.400 15.900 97.800 20.200 ;
        RECT 102.200 17.900 102.600 20.200 ;
        RECT 103.800 18.100 104.200 20.200 ;
        RECT 105.400 17.900 105.800 20.200 ;
        RECT 107.000 17.900 107.400 20.200 ;
        RECT 108.100 17.900 108.500 20.200 ;
        RECT 110.200 15.900 110.600 20.200 ;
        RECT 111.000 17.900 111.400 20.200 ;
        RECT 112.600 16.100 113.000 20.200 ;
        RECT 115.000 16.900 115.400 20.200 ;
        RECT 122.200 16.500 122.600 20.200 ;
        RECT 123.800 15.900 124.200 20.200 ;
        RECT 126.200 17.900 126.600 20.200 ;
        RECT 127.800 18.100 128.200 20.200 ;
        RECT 130.200 16.600 130.700 20.200 ;
        RECT 133.300 19.900 133.700 20.200 ;
        RECT 133.300 16.600 133.800 19.900 ;
        RECT 135.800 16.000 136.200 20.200 ;
        RECT 138.600 17.900 139.000 20.200 ;
        RECT 140.200 17.900 140.600 20.200 ;
        RECT 143.000 15.900 143.400 20.200 ;
        RECT 145.400 16.500 145.800 20.200 ;
        RECT 147.000 15.900 147.400 20.200 ;
        RECT 149.100 17.900 149.500 20.200 ;
        RECT 1.400 1.100 1.900 4.400 ;
        RECT 1.500 0.800 1.900 1.100 ;
        RECT 4.500 0.800 5.000 4.400 ;
        RECT 6.200 0.800 6.600 3.100 ;
        RECT 7.800 0.800 8.200 3.100 ;
        RECT 8.900 0.800 9.300 3.100 ;
        RECT 11.000 0.800 11.400 5.100 ;
        RECT 12.600 0.800 13.100 4.400 ;
        RECT 15.700 1.100 16.200 4.400 ;
        RECT 15.700 0.800 16.100 1.100 ;
        RECT 17.700 0.800 18.100 3.100 ;
        RECT 19.800 0.800 20.200 5.100 ;
        RECT 21.400 0.800 21.800 3.100 ;
        RECT 23.000 1.100 23.500 4.400 ;
        RECT 23.100 0.800 23.500 1.100 ;
        RECT 26.100 0.800 26.600 4.400 ;
        RECT 28.100 0.800 28.500 3.100 ;
        RECT 30.200 0.800 30.600 5.100 ;
        RECT 32.600 0.800 33.000 5.100 ;
        RECT 34.200 0.800 34.600 3.100 ;
        RECT 35.800 1.100 36.300 4.400 ;
        RECT 35.900 0.800 36.300 1.100 ;
        RECT 38.900 0.800 39.400 4.400 ;
        RECT 41.400 0.800 41.800 5.000 ;
        RECT 44.200 0.800 44.600 3.100 ;
        RECT 45.800 0.800 46.200 3.100 ;
        RECT 48.600 0.800 49.000 5.100 ;
        RECT 52.600 0.800 53.000 5.000 ;
        RECT 55.400 0.800 55.800 3.100 ;
        RECT 57.000 0.800 57.400 3.100 ;
        RECT 59.800 0.800 60.200 5.100 ;
        RECT 62.200 0.800 62.600 4.500 ;
        RECT 64.600 0.800 65.000 5.100 ;
        RECT 67.400 0.800 67.800 3.100 ;
        RECT 69.000 0.800 69.400 3.100 ;
        RECT 71.800 0.800 72.200 5.000 ;
        RECT 74.200 0.800 74.600 4.500 ;
        RECT 76.600 0.800 77.000 5.100 ;
        RECT 79.400 0.800 79.800 3.100 ;
        RECT 81.000 0.800 81.400 3.100 ;
        RECT 83.800 0.800 84.200 5.000 ;
        RECT 86.200 0.800 86.600 5.000 ;
        RECT 89.000 0.800 89.400 3.100 ;
        RECT 90.600 0.800 91.000 3.100 ;
        RECT 93.400 0.800 93.800 5.100 ;
        RECT 95.800 0.800 96.200 4.500 ;
        RECT 99.800 0.800 100.200 5.000 ;
        RECT 102.600 0.800 103.000 3.100 ;
        RECT 104.200 0.800 104.600 3.100 ;
        RECT 107.000 0.800 107.400 5.100 ;
        RECT 109.400 0.800 109.800 4.500 ;
        RECT 111.800 0.800 112.200 5.000 ;
        RECT 114.600 0.800 115.000 3.100 ;
        RECT 116.200 0.800 116.600 3.100 ;
        RECT 119.000 0.800 119.400 5.100 ;
        RECT 121.400 0.800 121.800 4.500 ;
        RECT 123.800 0.800 124.200 5.000 ;
        RECT 126.600 0.800 127.000 3.100 ;
        RECT 128.200 0.800 128.600 3.100 ;
        RECT 131.000 0.800 131.400 5.100 ;
        RECT 133.400 0.800 133.800 4.500 ;
        RECT 135.800 0.800 136.200 5.000 ;
        RECT 138.600 0.800 139.000 3.100 ;
        RECT 140.200 0.800 140.600 3.100 ;
        RECT 143.000 0.800 143.400 5.100 ;
        RECT 145.400 0.800 145.800 4.500 ;
        RECT 147.000 0.800 147.400 3.100 ;
        RECT 148.600 0.800 149.000 3.100 ;
        RECT 0.200 0.200 151.800 0.800 ;
      LAYER via1 ;
        RECT 49.000 120.300 49.400 120.700 ;
        RECT 49.700 120.300 50.100 120.700 ;
        RECT 49.000 100.300 49.400 100.700 ;
        RECT 49.700 100.300 50.100 100.700 ;
        RECT 49.000 80.300 49.400 80.700 ;
        RECT 49.700 80.300 50.100 80.700 ;
        RECT 49.000 60.300 49.400 60.700 ;
        RECT 49.700 60.300 50.100 60.700 ;
        RECT 49.000 40.300 49.400 40.700 ;
        RECT 49.700 40.300 50.100 40.700 ;
        RECT 49.000 20.300 49.400 20.700 ;
        RECT 49.700 20.300 50.100 20.700 ;
        RECT 49.000 0.300 49.400 0.700 ;
        RECT 49.700 0.300 50.100 0.700 ;
      LAYER metal2 ;
        RECT 48.800 120.300 50.400 120.700 ;
        RECT 48.800 100.300 50.400 100.700 ;
        RECT 48.800 80.300 50.400 80.700 ;
        RECT 48.800 60.300 50.400 60.700 ;
        RECT 48.800 40.300 50.400 40.700 ;
        RECT 48.800 20.300 50.400 20.700 ;
        RECT 48.800 0.300 50.400 0.700 ;
      LAYER via2 ;
        RECT 49.000 120.300 49.400 120.700 ;
        RECT 49.700 120.300 50.100 120.700 ;
        RECT 49.000 100.300 49.400 100.700 ;
        RECT 49.700 100.300 50.100 100.700 ;
        RECT 49.000 80.300 49.400 80.700 ;
        RECT 49.700 80.300 50.100 80.700 ;
        RECT 49.000 60.300 49.400 60.700 ;
        RECT 49.700 60.300 50.100 60.700 ;
        RECT 49.000 40.300 49.400 40.700 ;
        RECT 49.700 40.300 50.100 40.700 ;
        RECT 49.000 20.300 49.400 20.700 ;
        RECT 49.700 20.300 50.100 20.700 ;
        RECT 49.000 0.300 49.400 0.700 ;
        RECT 49.700 0.300 50.100 0.700 ;
      LAYER metal3 ;
        RECT 48.800 120.300 50.400 120.700 ;
        RECT 48.800 100.300 50.400 100.700 ;
        RECT 48.800 80.300 50.400 80.700 ;
        RECT 48.800 60.300 50.400 60.700 ;
        RECT 48.800 40.300 50.400 40.700 ;
        RECT 48.800 20.300 50.400 20.700 ;
        RECT 48.800 0.300 50.400 0.700 ;
      LAYER via3 ;
        RECT 49.000 120.300 49.400 120.700 ;
        RECT 49.800 120.300 50.200 120.700 ;
        RECT 49.000 100.300 49.400 100.700 ;
        RECT 49.800 100.300 50.200 100.700 ;
        RECT 49.000 80.300 49.400 80.700 ;
        RECT 49.800 80.300 50.200 80.700 ;
        RECT 49.000 60.300 49.400 60.700 ;
        RECT 49.800 60.300 50.200 60.700 ;
        RECT 49.000 40.300 49.400 40.700 ;
        RECT 49.800 40.300 50.200 40.700 ;
        RECT 49.000 20.300 49.400 20.700 ;
        RECT 49.800 20.300 50.200 20.700 ;
        RECT 49.000 0.300 49.400 0.700 ;
        RECT 49.800 0.300 50.200 0.700 ;
      LAYER metal4 ;
        RECT 48.800 120.300 50.400 120.700 ;
        RECT 48.800 100.300 50.400 100.700 ;
        RECT 48.800 80.300 50.400 80.700 ;
        RECT 48.800 60.300 50.400 60.700 ;
        RECT 48.800 40.300 50.400 40.700 ;
        RECT 48.800 20.300 50.400 20.700 ;
        RECT 48.800 0.300 50.400 0.700 ;
      LAYER via4 ;
        RECT 49.000 120.300 49.400 120.700 ;
        RECT 49.700 120.300 50.100 120.700 ;
        RECT 49.000 100.300 49.400 100.700 ;
        RECT 49.700 100.300 50.100 100.700 ;
        RECT 49.000 80.300 49.400 80.700 ;
        RECT 49.700 80.300 50.100 80.700 ;
        RECT 49.000 60.300 49.400 60.700 ;
        RECT 49.700 60.300 50.100 60.700 ;
        RECT 49.000 40.300 49.400 40.700 ;
        RECT 49.700 40.300 50.100 40.700 ;
        RECT 49.000 20.300 49.400 20.700 ;
        RECT 49.700 20.300 50.100 20.700 ;
        RECT 49.000 0.300 49.400 0.700 ;
        RECT 49.700 0.300 50.100 0.700 ;
      LAYER metal5 ;
        RECT 48.800 120.200 50.400 120.700 ;
        RECT 48.800 100.200 50.400 100.700 ;
        RECT 48.800 80.200 50.400 80.700 ;
        RECT 48.800 60.200 50.400 60.700 ;
        RECT 48.800 40.200 50.400 40.700 ;
        RECT 48.800 20.200 50.400 20.700 ;
        RECT 48.800 0.200 50.400 0.700 ;
      LAYER via5 ;
        RECT 49.800 120.200 50.300 120.700 ;
        RECT 49.800 100.200 50.300 100.700 ;
        RECT 49.800 80.200 50.300 80.700 ;
        RECT 49.800 60.200 50.300 60.700 ;
        RECT 49.800 40.200 50.300 40.700 ;
        RECT 49.800 20.200 50.300 20.700 ;
        RECT 49.800 0.200 50.300 0.700 ;
      LAYER metal6 ;
        RECT 48.800 -3.000 50.400 133.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 130.200 151.800 130.800 ;
        RECT 0.600 128.900 1.000 130.200 ;
        RECT 2.200 128.900 2.600 130.200 ;
        RECT 4.300 128.000 4.700 130.200 ;
        RECT 6.200 128.900 6.600 130.200 ;
        RECT 7.800 128.900 8.200 130.200 ;
        RECT 8.600 128.900 9.000 130.200 ;
        RECT 10.700 127.900 11.100 130.200 ;
        RECT 12.600 128.200 13.100 130.200 ;
        RECT 15.700 129.900 16.100 130.200 ;
        RECT 15.700 128.200 16.200 129.900 ;
        RECT 19.000 128.300 19.400 130.200 ;
        RECT 21.400 128.900 21.800 130.200 ;
        RECT 23.000 128.900 23.400 130.200 ;
        RECT 24.600 128.200 25.100 130.200 ;
        RECT 27.700 129.900 28.100 130.200 ;
        RECT 27.700 128.200 28.200 129.900 ;
        RECT 31.000 127.900 31.400 130.200 ;
        RECT 32.600 127.900 33.000 130.200 ;
        RECT 35.300 128.900 35.800 130.200 ;
        RECT 37.000 128.900 37.400 130.200 ;
        RECT 39.800 128.000 40.200 130.200 ;
        RECT 41.400 128.900 41.800 130.200 ;
        RECT 43.000 128.900 43.400 130.200 ;
        RECT 44.900 128.000 45.300 130.200 ;
        RECT 47.000 128.900 47.400 130.200 ;
        RECT 48.600 128.900 49.000 130.200 ;
        RECT 51.000 127.900 51.400 130.200 ;
        RECT 53.400 128.900 53.800 130.200 ;
        RECT 55.800 128.200 56.300 130.200 ;
        RECT 58.900 129.900 59.300 130.200 ;
        RECT 58.900 128.200 59.400 129.900 ;
        RECT 61.400 127.900 61.800 130.200 ;
        RECT 64.100 128.900 64.600 130.200 ;
        RECT 65.800 128.900 66.200 130.200 ;
        RECT 68.600 128.000 69.000 130.200 ;
        RECT 71.000 128.200 71.500 130.200 ;
        RECT 74.100 129.900 74.500 130.200 ;
        RECT 76.700 129.900 77.100 130.200 ;
        RECT 74.100 128.200 74.600 129.900 ;
        RECT 76.600 128.200 77.100 129.900 ;
        RECT 79.700 128.200 80.200 130.200 ;
        RECT 81.400 127.900 81.800 130.200 ;
        RECT 83.800 128.200 84.300 130.200 ;
        RECT 86.900 129.900 87.300 130.200 ;
        RECT 86.900 128.200 87.400 129.900 ;
        RECT 88.600 126.900 89.000 130.200 ;
        RECT 93.400 128.300 93.800 130.200 ;
        RECT 97.400 126.900 97.800 130.200 ;
        RECT 99.800 128.300 100.200 130.200 ;
        RECT 106.200 129.100 106.600 130.200 ;
        RECT 107.800 128.900 108.200 130.200 ;
        RECT 110.200 128.300 110.600 130.200 ;
        RECT 113.400 128.200 113.900 130.200 ;
        RECT 116.500 129.900 116.900 130.200 ;
        RECT 116.500 128.200 117.000 129.900 ;
        RECT 118.500 127.900 118.900 130.200 ;
        RECT 120.600 128.900 121.000 130.200 ;
        RECT 121.400 128.900 121.800 130.200 ;
        RECT 123.000 126.900 123.400 130.200 ;
        RECT 127.000 128.200 127.500 130.200 ;
        RECT 130.100 129.900 130.500 130.200 ;
        RECT 130.100 128.200 130.600 129.900 ;
        RECT 131.800 126.900 132.200 130.200 ;
        RECT 135.000 128.900 135.400 130.200 ;
        RECT 137.100 127.900 137.500 130.200 ;
        RECT 139.000 128.300 139.400 130.200 ;
        RECT 142.200 128.200 142.700 130.200 ;
        RECT 145.300 129.900 145.700 130.200 ;
        RECT 145.300 128.200 145.800 129.900 ;
        RECT 147.000 128.900 147.400 130.200 ;
        RECT 148.600 128.900 149.000 130.200 ;
        RECT 0.600 110.800 1.000 113.100 ;
        RECT 3.800 110.800 4.300 112.800 ;
        RECT 6.900 111.100 7.400 112.800 ;
        RECT 6.900 110.800 7.300 111.100 ;
        RECT 8.600 110.800 9.000 112.100 ;
        RECT 10.200 110.800 10.600 112.100 ;
        RECT 11.800 110.800 12.300 112.800 ;
        RECT 14.900 111.100 15.400 112.800 ;
        RECT 14.900 110.800 15.300 111.100 ;
        RECT 16.600 110.800 17.000 112.100 ;
        RECT 19.000 110.800 19.400 112.700 ;
        RECT 23.000 110.800 23.400 113.100 ;
        RECT 24.600 110.800 25.100 112.800 ;
        RECT 27.700 111.100 28.200 112.800 ;
        RECT 27.700 110.800 28.100 111.100 ;
        RECT 30.200 110.800 30.600 113.100 ;
        RECT 32.900 110.800 33.400 112.100 ;
        RECT 34.600 110.800 35.000 112.100 ;
        RECT 37.400 110.800 37.800 113.000 ;
        RECT 39.000 110.800 39.400 112.100 ;
        RECT 40.600 110.800 41.000 112.100 ;
        RECT 41.400 110.800 41.800 112.100 ;
        RECT 43.000 110.800 43.400 112.100 ;
        RECT 44.600 110.800 45.000 112.100 ;
        RECT 46.200 110.800 46.600 112.100 ;
        RECT 47.000 110.800 47.400 112.100 ;
        RECT 48.600 110.800 49.000 112.100 ;
        RECT 51.800 110.800 52.200 112.700 ;
        RECT 54.200 110.800 54.600 113.100 ;
        RECT 56.600 110.800 57.000 112.100 ;
        RECT 58.200 110.800 58.600 112.100 ;
        RECT 59.000 110.800 59.400 112.100 ;
        RECT 60.600 110.800 61.000 112.100 ;
        RECT 62.200 110.800 62.600 112.100 ;
        RECT 63.800 110.800 64.200 113.100 ;
        RECT 66.500 110.800 67.000 112.100 ;
        RECT 68.200 110.800 68.600 112.100 ;
        RECT 71.000 110.800 71.400 113.000 ;
        RECT 73.400 111.100 73.900 112.800 ;
        RECT 73.500 110.800 73.900 111.100 ;
        RECT 76.500 110.800 77.000 112.800 ;
        RECT 81.400 110.800 81.800 111.900 ;
        RECT 83.000 110.800 83.400 112.100 ;
        RECT 85.400 110.800 85.800 112.700 ;
        RECT 88.600 110.800 89.000 112.100 ;
        RECT 89.400 110.800 89.800 114.100 ;
        RECT 92.600 110.800 93.000 112.100 ;
        RECT 96.600 110.800 97.000 114.100 ;
        RECT 97.400 110.800 97.800 112.100 ;
        RECT 99.500 110.800 99.900 113.100 ;
        RECT 102.500 110.800 102.900 113.100 ;
        RECT 104.600 110.800 105.000 112.100 ;
        RECT 106.200 110.800 106.600 112.100 ;
        RECT 107.800 110.800 108.200 111.900 ;
        RECT 112.600 110.800 113.000 112.700 ;
        RECT 115.800 111.100 116.300 112.800 ;
        RECT 115.900 110.800 116.300 111.100 ;
        RECT 118.900 110.800 119.400 112.800 ;
        RECT 120.600 110.800 121.000 114.100 ;
        RECT 126.200 110.800 126.600 114.100 ;
        RECT 127.300 110.800 127.700 113.100 ;
        RECT 129.400 110.800 129.800 112.100 ;
        RECT 131.000 110.800 131.500 112.800 ;
        RECT 134.100 111.100 134.600 112.800 ;
        RECT 134.100 110.800 134.500 111.100 ;
        RECT 138.200 110.800 138.600 114.100 ;
        RECT 139.300 110.800 139.700 113.100 ;
        RECT 141.400 110.800 141.800 112.100 ;
        RECT 144.600 110.800 145.000 114.100 ;
        RECT 146.200 110.800 146.600 112.100 ;
        RECT 147.000 110.800 147.400 112.100 ;
        RECT 149.100 110.800 149.500 113.100 ;
        RECT 0.200 110.200 151.800 110.800 ;
        RECT 0.600 108.900 1.000 110.200 ;
        RECT 2.200 108.900 2.600 110.200 ;
        RECT 3.000 108.900 3.400 110.200 ;
        RECT 4.600 108.900 5.000 110.200 ;
        RECT 6.200 108.900 6.600 110.200 ;
        RECT 7.800 108.900 8.200 110.200 ;
        RECT 8.600 107.900 9.000 110.200 ;
        RECT 11.800 107.900 12.200 110.200 ;
        RECT 14.500 108.900 15.000 110.200 ;
        RECT 16.200 108.900 16.600 110.200 ;
        RECT 19.000 108.000 19.400 110.200 ;
        RECT 21.400 107.900 21.800 110.200 ;
        RECT 24.100 108.900 24.600 110.200 ;
        RECT 25.800 108.900 26.200 110.200 ;
        RECT 28.600 108.000 29.000 110.200 ;
        RECT 31.100 109.900 31.500 110.200 ;
        RECT 31.000 108.200 31.500 109.900 ;
        RECT 34.100 108.200 34.600 110.200 ;
        RECT 35.800 107.900 36.200 110.200 ;
        RECT 39.000 108.200 39.500 110.200 ;
        RECT 42.100 109.900 42.500 110.200 ;
        RECT 42.100 108.200 42.600 109.900 ;
        RECT 43.800 108.900 44.200 110.200 ;
        RECT 47.000 108.300 47.400 110.200 ;
        RECT 51.000 108.200 51.500 110.200 ;
        RECT 54.100 109.900 54.500 110.200 ;
        RECT 54.100 108.200 54.600 109.900 ;
        RECT 56.600 107.900 57.000 110.200 ;
        RECT 59.300 108.900 59.800 110.200 ;
        RECT 61.000 108.900 61.400 110.200 ;
        RECT 63.800 108.000 64.200 110.200 ;
        RECT 66.200 107.900 66.600 110.200 ;
        RECT 68.900 108.900 69.400 110.200 ;
        RECT 70.600 108.900 71.000 110.200 ;
        RECT 73.400 108.000 73.800 110.200 ;
        RECT 75.900 109.900 76.300 110.200 ;
        RECT 75.800 108.200 76.300 109.900 ;
        RECT 78.900 108.200 79.400 110.200 ;
        RECT 80.600 107.900 81.000 110.200 ;
        RECT 83.300 107.900 83.700 110.200 ;
        RECT 85.400 108.900 85.800 110.200 ;
        RECT 88.600 106.900 89.000 110.200 ;
        RECT 91.800 106.900 92.200 110.200 ;
        RECT 92.600 108.900 93.000 110.200 ;
        RECT 94.700 107.900 95.100 110.200 ;
        RECT 96.100 107.900 96.500 110.200 ;
        RECT 98.200 108.900 98.600 110.200 ;
        RECT 99.000 107.900 99.400 110.200 ;
        RECT 105.400 106.900 105.800 110.200 ;
        RECT 108.600 106.900 109.000 110.200 ;
        RECT 109.400 108.900 109.800 110.200 ;
        RECT 112.600 108.300 113.000 110.200 ;
        RECT 115.000 108.300 115.400 110.200 ;
        RECT 119.800 106.900 120.200 110.200 ;
        RECT 120.900 107.900 121.300 110.200 ;
        RECT 123.000 108.900 123.400 110.200 ;
        RECT 124.600 108.300 125.000 110.200 ;
        RECT 129.400 106.900 129.800 110.200 ;
        RECT 130.500 107.900 130.900 110.200 ;
        RECT 132.600 108.900 133.000 110.200 ;
        RECT 133.400 108.900 133.800 110.200 ;
        RECT 135.500 107.900 135.900 110.200 ;
        RECT 137.400 108.200 137.900 110.200 ;
        RECT 140.500 109.900 140.900 110.200 ;
        RECT 140.500 108.200 141.000 109.900 ;
        RECT 143.000 108.300 143.400 110.200 ;
        RECT 147.800 106.900 148.200 110.200 ;
        RECT 148.900 107.900 149.300 110.200 ;
        RECT 151.000 108.900 151.400 110.200 ;
        RECT 0.600 90.800 1.000 92.100 ;
        RECT 3.800 90.800 4.200 93.100 ;
        RECT 4.600 90.800 5.000 92.100 ;
        RECT 6.200 90.800 6.600 92.100 ;
        RECT 7.000 90.800 7.400 92.100 ;
        RECT 9.900 90.800 10.300 93.000 ;
        RECT 12.600 90.800 13.100 92.800 ;
        RECT 15.700 91.100 16.200 92.800 ;
        RECT 15.700 90.800 16.100 91.100 ;
        RECT 18.200 90.800 18.600 93.100 ;
        RECT 20.900 90.800 21.400 92.100 ;
        RECT 22.600 90.800 23.000 92.100 ;
        RECT 25.400 90.800 25.800 93.000 ;
        RECT 27.800 90.800 28.200 93.100 ;
        RECT 30.500 90.800 31.000 92.100 ;
        RECT 32.200 90.800 32.600 92.100 ;
        RECT 35.000 90.800 35.400 93.000 ;
        RECT 36.600 90.800 37.000 92.100 ;
        RECT 38.200 90.800 38.600 92.100 ;
        RECT 39.000 90.800 39.400 93.100 ;
        RECT 42.200 90.800 42.600 93.100 ;
        RECT 44.900 90.800 45.400 92.100 ;
        RECT 46.600 90.800 47.000 92.100 ;
        RECT 49.400 90.800 49.800 93.000 ;
        RECT 52.600 90.800 53.000 92.100 ;
        RECT 54.200 90.800 54.600 92.100 ;
        RECT 55.800 90.800 56.200 92.100 ;
        RECT 56.600 90.800 57.000 92.100 ;
        RECT 58.700 90.800 59.100 93.100 ;
        RECT 59.800 90.800 60.200 94.100 ;
        RECT 63.000 90.800 63.400 92.100 ;
        RECT 64.600 90.800 65.000 92.100 ;
        RECT 66.200 90.800 66.600 92.700 ;
        RECT 70.200 90.800 70.600 92.700 ;
        RECT 73.400 90.800 73.800 92.700 ;
        RECT 76.600 90.800 77.000 92.100 ;
        RECT 79.000 90.800 79.400 92.700 ;
        RECT 81.400 90.800 81.800 92.700 ;
        RECT 83.800 90.800 84.200 93.100 ;
        RECT 86.200 90.800 86.600 93.100 ;
        RECT 90.200 90.800 90.600 93.100 ;
        RECT 91.000 90.800 91.400 94.100 ;
        RECT 94.200 90.800 94.600 93.100 ;
        RECT 96.600 90.800 97.000 93.100 ;
        RECT 101.400 90.800 101.800 92.700 ;
        RECT 104.800 90.800 105.200 93.100 ;
        RECT 107.800 90.800 108.200 93.100 ;
        RECT 108.600 90.800 109.000 93.100 ;
        RECT 111.000 90.800 111.400 94.100 ;
        RECT 114.500 90.800 114.900 93.100 ;
        RECT 116.600 90.800 117.000 92.100 ;
        RECT 117.400 90.800 117.800 92.100 ;
        RECT 119.000 90.800 119.400 92.100 ;
        RECT 120.600 90.800 121.000 92.700 ;
        RECT 123.000 90.800 123.400 94.100 ;
        RECT 128.600 90.800 129.000 94.100 ;
        RECT 131.800 90.800 132.200 94.100 ;
        RECT 135.000 90.800 135.400 94.100 ;
        RECT 135.800 90.800 136.200 94.100 ;
        RECT 139.000 90.800 139.400 94.100 ;
        RECT 142.500 90.800 142.900 93.100 ;
        RECT 144.600 90.800 145.000 92.100 ;
        RECT 145.400 90.800 145.800 93.100 ;
        RECT 150.200 90.800 150.600 94.100 ;
        RECT 0.200 90.200 151.800 90.800 ;
        RECT 0.600 88.900 1.000 90.200 ;
        RECT 2.200 87.900 2.600 90.200 ;
        RECT 4.600 88.900 5.000 90.200 ;
        RECT 6.200 88.100 6.600 90.200 ;
        RECT 9.100 88.000 9.500 90.200 ;
        RECT 12.600 88.300 13.000 90.200 ;
        RECT 14.200 88.900 14.600 90.200 ;
        RECT 15.800 88.900 16.200 90.200 ;
        RECT 17.900 87.900 18.300 90.200 ;
        RECT 19.000 88.900 19.400 90.200 ;
        RECT 20.600 88.900 21.000 90.200 ;
        RECT 21.400 87.900 21.800 90.200 ;
        RECT 23.800 88.200 24.300 90.200 ;
        RECT 26.900 89.900 27.300 90.200 ;
        RECT 26.900 88.200 27.400 89.900 ;
        RECT 29.400 87.900 29.800 90.200 ;
        RECT 32.100 88.900 32.600 90.200 ;
        RECT 33.800 88.900 34.200 90.200 ;
        RECT 36.600 88.000 37.000 90.200 ;
        RECT 39.000 87.900 39.400 90.200 ;
        RECT 41.700 88.900 42.200 90.200 ;
        RECT 43.400 88.900 43.800 90.200 ;
        RECT 46.200 88.000 46.600 90.200 ;
        RECT 50.200 87.900 50.600 90.200 ;
        RECT 52.900 88.900 53.400 90.200 ;
        RECT 54.600 88.900 55.000 90.200 ;
        RECT 57.400 88.000 57.800 90.200 ;
        RECT 59.000 88.900 59.400 90.200 ;
        RECT 61.900 88.000 62.300 90.200 ;
        RECT 63.800 87.900 64.200 90.200 ;
        RECT 66.200 87.900 66.600 90.200 ;
        RECT 70.200 87.900 70.600 90.200 ;
        RECT 71.000 87.900 71.400 90.200 ;
        RECT 74.000 87.900 74.400 90.200 ;
        RECT 75.000 87.900 75.400 90.200 ;
        RECT 77.400 87.900 77.800 90.200 ;
        RECT 79.800 88.900 80.200 90.200 ;
        RECT 81.900 87.900 82.300 90.200 ;
        RECT 83.800 88.900 84.200 90.200 ;
        RECT 84.900 87.900 85.300 90.200 ;
        RECT 87.000 88.900 87.400 90.200 ;
        RECT 87.800 87.900 88.200 90.200 ;
        RECT 90.200 88.900 90.600 90.200 ;
        RECT 92.600 88.300 93.000 90.200 ;
        RECT 95.000 87.900 95.400 90.200 ;
        RECT 98.000 87.900 98.400 90.200 ;
        RECT 99.000 87.900 99.400 90.200 ;
        RECT 104.600 87.900 105.000 90.200 ;
        RECT 105.400 86.900 105.800 90.200 ;
        RECT 108.900 87.900 109.300 90.200 ;
        RECT 111.000 88.900 111.400 90.200 ;
        RECT 111.800 86.900 112.200 90.200 ;
        RECT 115.300 87.900 115.700 90.200 ;
        RECT 117.400 88.900 117.800 90.200 ;
        RECT 119.000 88.300 119.400 90.200 ;
        RECT 122.200 88.900 122.600 90.200 ;
        RECT 123.800 88.900 124.200 90.200 ;
        RECT 126.200 88.300 126.600 90.200 ;
        RECT 128.600 88.300 129.000 90.200 ;
        RECT 131.000 88.900 131.400 90.200 ;
        RECT 133.100 87.900 133.500 90.200 ;
        RECT 136.600 86.900 137.000 90.200 ;
        RECT 139.800 86.900 140.200 90.200 ;
        RECT 140.900 87.900 141.300 90.200 ;
        RECT 143.000 88.900 143.400 90.200 ;
        RECT 143.800 86.900 144.200 90.200 ;
        RECT 147.000 86.900 147.400 90.200 ;
        RECT 0.600 70.800 1.000 72.100 ;
        RECT 2.200 70.800 2.600 72.100 ;
        RECT 3.800 70.800 4.200 72.100 ;
        RECT 5.400 70.800 5.800 72.100 ;
        RECT 7.000 71.100 7.500 72.800 ;
        RECT 7.100 70.800 7.500 71.100 ;
        RECT 10.100 70.800 10.600 72.800 ;
        RECT 11.800 70.800 12.200 72.100 ;
        RECT 14.200 70.800 14.600 72.700 ;
        RECT 16.600 70.800 17.000 72.100 ;
        RECT 18.700 70.800 19.100 73.100 ;
        RECT 20.600 70.800 21.000 73.100 ;
        RECT 23.300 70.800 23.800 72.100 ;
        RECT 25.000 70.800 25.400 72.100 ;
        RECT 27.800 70.800 28.200 73.000 ;
        RECT 30.200 70.800 30.600 73.100 ;
        RECT 32.900 70.800 33.400 72.100 ;
        RECT 34.600 70.800 35.000 72.100 ;
        RECT 37.400 70.800 37.800 73.000 ;
        RECT 39.800 70.800 40.200 73.100 ;
        RECT 42.500 70.800 43.000 72.100 ;
        RECT 44.200 70.800 44.600 72.100 ;
        RECT 47.000 70.800 47.400 73.000 ;
        RECT 51.000 70.800 51.400 73.100 ;
        RECT 53.700 70.800 54.200 72.100 ;
        RECT 55.400 70.800 55.800 72.100 ;
        RECT 58.200 70.800 58.600 73.000 ;
        RECT 59.800 70.800 60.200 73.100 ;
        RECT 64.600 70.800 65.000 74.100 ;
        RECT 65.400 70.800 65.800 72.100 ;
        RECT 67.500 70.800 67.900 73.100 ;
        RECT 68.600 70.800 69.000 73.100 ;
        RECT 71.000 70.800 71.400 72.100 ;
        RECT 73.100 70.800 73.500 73.100 ;
        RECT 75.000 70.800 75.400 73.100 ;
        RECT 76.600 70.800 77.000 73.100 ;
        RECT 78.200 70.800 78.600 73.100 ;
        RECT 79.800 70.800 80.200 73.100 ;
        RECT 81.400 70.800 81.800 73.100 ;
        RECT 83.000 70.800 83.400 73.100 ;
        RECT 83.800 70.800 84.200 73.100 ;
        RECT 86.400 70.800 86.800 73.100 ;
        RECT 89.400 70.800 89.800 73.100 ;
        RECT 90.200 70.800 90.600 73.100 ;
        RECT 92.600 70.800 93.000 73.100 ;
        RECT 95.600 70.800 96.000 73.100 ;
        RECT 96.900 70.800 97.300 73.100 ;
        RECT 99.000 70.800 99.400 72.100 ;
        RECT 101.700 70.800 102.100 73.100 ;
        RECT 103.800 70.800 104.200 72.100 ;
        RECT 104.600 70.800 105.000 73.100 ;
        RECT 107.000 70.800 107.400 72.100 ;
        RECT 108.600 70.800 109.000 72.100 ;
        RECT 109.400 70.800 109.800 73.100 ;
        RECT 114.200 70.800 114.600 74.100 ;
        RECT 117.400 70.800 117.800 74.100 ;
        RECT 119.000 70.800 119.400 73.100 ;
        RECT 119.800 70.800 120.200 74.100 ;
        RECT 123.300 70.800 123.700 73.100 ;
        RECT 125.400 70.800 125.800 72.100 ;
        RECT 126.200 70.800 126.600 74.100 ;
        RECT 130.200 70.800 130.600 72.700 ;
        RECT 133.400 71.100 133.900 72.800 ;
        RECT 133.500 70.800 133.900 71.100 ;
        RECT 136.500 70.800 137.000 72.800 ;
        RECT 138.200 70.800 138.600 74.100 ;
        RECT 141.400 70.800 141.800 74.100 ;
        RECT 147.000 70.800 147.400 74.100 ;
        RECT 148.100 70.800 148.500 73.100 ;
        RECT 150.200 70.800 150.600 72.100 ;
        RECT 0.200 70.200 151.800 70.800 ;
        RECT 0.600 68.900 1.000 70.200 ;
        RECT 2.200 68.900 2.600 70.200 ;
        RECT 3.800 68.200 4.300 70.200 ;
        RECT 6.900 69.900 7.300 70.200 ;
        RECT 6.900 68.200 7.400 69.900 ;
        RECT 8.600 68.900 9.000 70.200 ;
        RECT 10.500 67.900 10.900 70.200 ;
        RECT 12.600 68.900 13.000 70.200 ;
        RECT 13.400 68.900 13.800 70.200 ;
        RECT 15.000 68.900 15.400 70.200 ;
        RECT 17.400 67.900 17.800 70.200 ;
        RECT 19.000 68.200 19.500 70.200 ;
        RECT 22.100 69.900 22.500 70.200 ;
        RECT 22.100 68.200 22.600 69.900 ;
        RECT 24.600 68.200 25.100 70.200 ;
        RECT 27.700 69.900 28.100 70.200 ;
        RECT 27.700 68.200 28.200 69.900 ;
        RECT 30.200 68.200 30.700 70.200 ;
        RECT 33.300 69.900 33.700 70.200 ;
        RECT 33.300 68.200 33.800 69.900 ;
        RECT 35.000 68.900 35.400 70.200 ;
        RECT 36.600 68.900 37.000 70.200 ;
        RECT 38.200 67.900 38.600 70.200 ;
        RECT 40.900 68.900 41.400 70.200 ;
        RECT 42.600 68.900 43.000 70.200 ;
        RECT 45.400 68.000 45.800 70.200 ;
        RECT 49.400 67.900 49.800 70.200 ;
        RECT 52.100 68.900 52.600 70.200 ;
        RECT 53.800 68.900 54.200 70.200 ;
        RECT 56.600 68.000 57.000 70.200 ;
        RECT 58.200 67.900 58.600 70.200 ;
        RECT 60.600 67.900 61.000 70.200 ;
        RECT 65.400 66.900 65.800 70.200 ;
        RECT 68.600 66.900 69.000 70.200 ;
        RECT 69.400 68.900 69.800 70.200 ;
        RECT 72.600 68.300 73.000 70.200 ;
        RECT 75.000 68.300 75.400 70.200 ;
        RECT 77.400 67.900 77.800 70.200 ;
        RECT 79.800 67.900 80.200 70.200 ;
        RECT 82.200 67.900 82.600 70.200 ;
        RECT 83.800 67.900 84.200 70.200 ;
        RECT 86.200 67.900 86.600 70.200 ;
        RECT 87.800 67.900 88.200 70.200 ;
        RECT 90.200 67.900 90.600 70.200 ;
        RECT 91.800 68.300 92.200 70.200 ;
        RECT 96.600 68.300 97.000 70.200 ;
        RECT 99.000 68.300 99.400 70.200 ;
        RECT 103.000 67.900 103.400 70.200 ;
        RECT 106.200 68.300 106.600 70.200 ;
        RECT 108.600 68.300 109.000 70.200 ;
        RECT 111.300 67.900 111.700 70.200 ;
        RECT 113.400 68.900 113.800 70.200 ;
        RECT 114.200 66.900 114.600 70.200 ;
        RECT 119.800 66.900 120.200 70.200 ;
        RECT 120.600 66.900 121.000 70.200 ;
        RECT 124.100 67.900 124.500 70.200 ;
        RECT 126.200 68.900 126.600 70.200 ;
        RECT 127.000 66.900 127.400 70.200 ;
        RECT 130.200 66.900 130.600 70.200 ;
        RECT 133.400 66.900 133.800 70.200 ;
        RECT 136.900 67.900 137.300 70.200 ;
        RECT 139.000 68.900 139.400 70.200 ;
        RECT 142.200 66.900 142.600 70.200 ;
        RECT 145.400 66.900 145.800 70.200 ;
        RECT 147.000 68.200 147.500 70.200 ;
        RECT 150.100 69.900 150.500 70.200 ;
        RECT 150.100 68.200 150.600 69.900 ;
        RECT 1.400 51.100 1.900 52.800 ;
        RECT 1.500 50.800 1.900 51.100 ;
        RECT 4.500 50.800 5.000 52.800 ;
        RECT 7.000 50.800 7.400 53.100 ;
        RECT 9.700 50.800 10.200 52.100 ;
        RECT 11.400 50.800 11.800 52.100 ;
        RECT 14.200 50.800 14.600 53.000 ;
        RECT 16.600 51.100 17.100 52.800 ;
        RECT 16.700 50.800 17.100 51.100 ;
        RECT 19.700 50.800 20.200 52.800 ;
        RECT 21.400 50.800 21.800 53.100 ;
        RECT 23.800 50.800 24.200 52.100 ;
        RECT 25.400 50.800 25.800 52.100 ;
        RECT 27.000 50.800 27.400 52.100 ;
        RECT 27.800 50.800 28.200 52.100 ;
        RECT 29.400 50.800 29.800 52.100 ;
        RECT 30.200 50.800 30.600 52.100 ;
        RECT 31.800 50.800 32.200 53.100 ;
        RECT 33.400 50.800 33.800 53.100 ;
        RECT 35.000 50.800 35.400 53.100 ;
        RECT 36.600 50.800 37.000 53.100 ;
        RECT 38.200 50.800 38.600 53.100 ;
        RECT 39.800 50.800 40.200 53.100 ;
        RECT 42.500 50.800 43.000 52.100 ;
        RECT 44.200 50.800 44.600 52.100 ;
        RECT 47.000 50.800 47.400 53.000 ;
        RECT 50.500 50.800 50.900 53.100 ;
        RECT 52.600 50.800 53.000 52.100 ;
        RECT 55.800 50.800 56.200 54.100 ;
        RECT 56.600 50.800 57.000 53.100 ;
        RECT 59.000 50.800 59.400 53.100 ;
        RECT 61.400 50.800 61.800 53.100 ;
        RECT 65.400 50.800 65.800 53.100 ;
        RECT 67.000 50.800 67.400 53.100 ;
        RECT 68.600 50.800 69.000 53.100 ;
        RECT 70.200 50.800 70.600 52.700 ;
        RECT 72.600 50.800 73.000 53.100 ;
        RECT 76.600 50.800 77.000 53.100 ;
        RECT 77.400 50.800 77.800 53.100 ;
        RECT 81.400 50.800 81.800 53.100 ;
        RECT 82.200 50.800 82.600 52.100 ;
        RECT 83.800 50.800 84.200 52.100 ;
        RECT 85.400 50.800 85.800 52.700 ;
        RECT 88.600 50.800 89.000 52.100 ;
        RECT 90.700 50.800 91.100 53.100 ;
        RECT 91.800 50.800 92.200 54.100 ;
        RECT 97.400 50.800 97.800 54.100 ;
        RECT 98.500 50.800 98.900 53.100 ;
        RECT 100.600 50.800 101.000 52.100 ;
        RECT 103.800 50.800 104.200 52.700 ;
        RECT 108.600 50.800 109.000 54.100 ;
        RECT 109.700 50.800 110.100 53.100 ;
        RECT 111.800 50.800 112.200 52.100 ;
        RECT 112.600 50.800 113.000 54.100 ;
        RECT 118.200 50.800 118.600 54.100 ;
        RECT 119.300 50.800 119.700 53.100 ;
        RECT 121.400 50.800 121.800 52.100 ;
        RECT 124.600 50.800 125.000 54.100 ;
        RECT 125.400 50.800 125.800 52.100 ;
        RECT 127.500 50.800 127.900 53.100 ;
        RECT 129.400 50.800 129.800 52.700 ;
        RECT 134.200 50.800 134.600 54.100 ;
        RECT 135.000 50.800 135.400 54.100 ;
        RECT 138.200 50.800 138.600 53.100 ;
        RECT 141.400 50.800 141.800 53.100 ;
        RECT 143.000 50.800 143.500 52.800 ;
        RECT 146.100 51.100 146.600 52.800 ;
        RECT 146.100 50.800 146.500 51.100 ;
        RECT 148.600 50.800 149.000 52.700 ;
        RECT 0.200 50.200 151.800 50.800 ;
        RECT 0.600 47.900 1.000 50.200 ;
        RECT 3.800 48.200 4.300 50.200 ;
        RECT 6.900 49.900 7.300 50.200 ;
        RECT 6.900 48.200 7.400 49.900 ;
        RECT 10.200 48.300 10.600 50.200 ;
        RECT 12.600 48.200 13.100 50.200 ;
        RECT 15.700 49.900 16.100 50.200 ;
        RECT 15.700 48.200 16.200 49.900 ;
        RECT 18.200 47.900 18.600 50.200 ;
        RECT 20.900 48.900 21.400 50.200 ;
        RECT 22.600 48.900 23.000 50.200 ;
        RECT 25.400 48.000 25.800 50.200 ;
        RECT 27.000 47.900 27.400 50.200 ;
        RECT 28.600 47.900 29.000 50.200 ;
        RECT 30.200 47.900 30.600 50.200 ;
        RECT 31.800 47.900 32.200 50.200 ;
        RECT 33.400 47.900 33.800 50.200 ;
        RECT 34.200 48.900 34.600 50.200 ;
        RECT 35.800 48.900 36.200 50.200 ;
        RECT 37.900 48.000 38.300 50.200 ;
        RECT 40.600 48.300 41.000 50.200 ;
        RECT 43.800 48.900 44.200 50.200 ;
        RECT 44.600 48.900 45.000 50.200 ;
        RECT 46.200 48.900 46.600 50.200 ;
        RECT 47.000 48.900 47.400 50.200 ;
        RECT 49.100 47.900 49.500 50.200 ;
        RECT 52.600 48.200 53.100 50.200 ;
        RECT 55.700 49.900 56.100 50.200 ;
        RECT 55.700 48.200 56.200 49.900 ;
        RECT 58.200 47.900 58.600 50.200 ;
        RECT 60.900 48.900 61.400 50.200 ;
        RECT 62.600 48.900 63.000 50.200 ;
        RECT 65.400 48.000 65.800 50.200 ;
        RECT 67.000 47.900 67.400 50.200 ;
        RECT 68.600 47.900 69.000 50.200 ;
        RECT 70.200 47.900 70.600 50.200 ;
        RECT 71.800 47.900 72.200 50.200 ;
        RECT 73.400 47.900 73.800 50.200 ;
        RECT 74.200 48.900 74.600 50.200 ;
        RECT 75.800 48.900 76.200 50.200 ;
        RECT 78.200 48.300 78.600 50.200 ;
        RECT 80.600 48.900 81.000 50.200 ;
        RECT 83.000 48.300 83.400 50.200 ;
        RECT 84.600 47.900 85.000 50.200 ;
        RECT 86.200 48.900 86.600 50.200 ;
        RECT 87.800 48.900 88.200 50.200 ;
        RECT 88.600 48.900 89.000 50.200 ;
        RECT 90.200 48.900 90.600 50.200 ;
        RECT 91.800 47.900 92.200 50.200 ;
        RECT 93.400 47.900 93.800 50.200 ;
        RECT 94.200 47.900 94.600 50.200 ;
        RECT 97.400 48.300 97.800 50.200 ;
        RECT 99.000 48.900 99.400 50.200 ;
        RECT 100.600 48.900 101.000 50.200 ;
        RECT 103.000 48.900 103.400 50.200 ;
        RECT 105.100 47.900 105.500 50.200 ;
        RECT 107.000 48.900 107.400 50.200 ;
        RECT 108.600 48.300 109.000 50.200 ;
        RECT 111.800 48.300 112.200 50.200 ;
        RECT 114.200 48.900 114.600 50.200 ;
        RECT 115.800 48.900 116.200 50.200 ;
        RECT 117.900 47.900 118.300 50.200 ;
        RECT 119.000 46.900 119.400 50.200 ;
        RECT 122.200 47.900 122.600 50.200 ;
        RECT 124.100 47.900 124.500 50.200 ;
        RECT 126.200 48.900 126.600 50.200 ;
        RECT 127.800 48.300 128.200 50.200 ;
        RECT 132.600 46.900 133.000 50.200 ;
        RECT 133.400 48.900 133.800 50.200 ;
        RECT 135.500 47.900 135.900 50.200 ;
        RECT 136.600 48.900 137.000 50.200 ;
        RECT 138.200 48.100 138.600 50.200 ;
        RECT 139.800 47.900 140.200 50.200 ;
        RECT 142.200 46.900 142.600 50.200 ;
        RECT 145.400 48.900 145.800 50.200 ;
        RECT 147.000 48.900 147.400 50.200 ;
        RECT 149.100 48.000 149.500 50.200 ;
        RECT 1.400 31.100 1.900 32.800 ;
        RECT 1.500 30.800 1.900 31.100 ;
        RECT 4.500 30.800 5.000 32.800 ;
        RECT 6.200 30.800 6.600 33.100 ;
        RECT 9.400 30.800 9.800 32.100 ;
        RECT 11.800 30.800 12.200 32.700 ;
        RECT 14.200 30.800 14.700 32.800 ;
        RECT 17.300 31.100 17.800 32.800 ;
        RECT 17.300 30.800 17.700 31.100 ;
        RECT 19.800 30.800 20.200 33.100 ;
        RECT 22.500 30.800 23.000 32.100 ;
        RECT 24.200 30.800 24.600 32.100 ;
        RECT 27.000 30.800 27.400 33.000 ;
        RECT 29.400 30.800 29.800 33.100 ;
        RECT 32.100 30.800 32.600 32.100 ;
        RECT 33.800 30.800 34.200 32.100 ;
        RECT 36.600 30.800 37.000 33.000 ;
        RECT 39.000 30.800 39.400 32.100 ;
        RECT 40.600 30.800 41.100 32.800 ;
        RECT 43.700 31.100 44.200 32.800 ;
        RECT 43.700 30.800 44.100 31.100 ;
        RECT 47.000 30.800 47.400 33.100 ;
        RECT 50.200 31.100 50.700 32.800 ;
        RECT 50.300 30.800 50.700 31.100 ;
        RECT 53.300 30.800 53.800 32.800 ;
        RECT 55.800 30.800 56.200 33.100 ;
        RECT 58.500 30.800 59.000 32.100 ;
        RECT 60.200 30.800 60.600 32.100 ;
        RECT 63.000 30.800 63.400 33.000 ;
        RECT 65.400 30.800 65.800 33.100 ;
        RECT 68.100 30.800 68.600 32.100 ;
        RECT 69.800 30.800 70.200 32.100 ;
        RECT 72.600 30.800 73.000 33.000 ;
        RECT 74.200 30.800 74.600 33.100 ;
        RECT 75.800 30.800 76.200 33.100 ;
        RECT 76.600 30.800 77.000 32.100 ;
        RECT 78.200 30.800 78.600 32.100 ;
        RECT 79.000 30.800 79.400 32.100 ;
        RECT 81.400 30.800 81.800 32.700 ;
        RECT 83.800 30.800 84.200 32.100 ;
        RECT 85.400 30.800 85.800 32.100 ;
        RECT 87.800 30.800 88.200 32.700 ;
        RECT 91.000 30.800 91.400 32.700 ;
        RECT 93.400 30.800 93.800 32.100 ;
        RECT 95.000 30.800 95.400 33.100 ;
        RECT 96.600 30.800 97.000 33.100 ;
        RECT 98.200 30.800 98.600 32.700 ;
        RECT 103.800 30.800 104.200 33.100 ;
        RECT 104.600 30.800 105.000 32.100 ;
        RECT 106.200 30.800 106.600 32.100 ;
        RECT 108.300 30.800 108.700 33.100 ;
        RECT 109.400 30.800 109.800 34.100 ;
        RECT 113.400 30.800 113.800 32.700 ;
        RECT 115.800 30.800 116.200 32.100 ;
        RECT 117.900 30.800 118.300 33.100 ;
        RECT 120.600 30.800 121.000 33.100 ;
        RECT 122.200 30.800 122.600 32.700 ;
        RECT 124.600 30.800 125.000 32.100 ;
        RECT 126.700 30.800 127.100 33.100 ;
        RECT 130.200 30.800 130.600 34.100 ;
        RECT 131.000 30.800 131.400 34.100 ;
        RECT 134.200 30.800 134.600 32.100 ;
        RECT 136.300 30.800 136.700 33.100 ;
        RECT 139.800 30.800 140.200 34.100 ;
        RECT 140.900 30.800 141.300 33.100 ;
        RECT 143.000 30.800 143.400 32.100 ;
        RECT 143.800 30.800 144.200 34.100 ;
        RECT 148.600 30.800 149.000 32.700 ;
        RECT 0.200 30.200 151.800 30.800 ;
        RECT 0.600 27.900 1.000 30.200 ;
        RECT 2.200 27.900 2.600 30.200 ;
        RECT 3.800 27.900 4.200 30.200 ;
        RECT 5.400 27.900 5.800 30.200 ;
        RECT 7.000 27.900 7.400 30.200 ;
        RECT 8.600 28.200 9.100 30.200 ;
        RECT 11.700 29.900 12.100 30.200 ;
        RECT 11.700 28.200 12.200 29.900 ;
        RECT 14.200 27.900 14.600 30.200 ;
        RECT 16.900 28.900 17.400 30.200 ;
        RECT 18.600 28.900 19.000 30.200 ;
        RECT 21.400 28.000 21.800 30.200 ;
        RECT 23.800 27.900 24.200 30.200 ;
        RECT 26.500 28.900 27.000 30.200 ;
        RECT 28.200 28.900 28.600 30.200 ;
        RECT 31.000 28.000 31.400 30.200 ;
        RECT 33.400 27.900 33.800 30.200 ;
        RECT 36.100 28.900 36.600 30.200 ;
        RECT 37.800 28.900 38.200 30.200 ;
        RECT 40.600 28.000 41.000 30.200 ;
        RECT 43.000 27.900 43.400 30.200 ;
        RECT 45.700 28.900 46.200 30.200 ;
        RECT 47.400 28.900 47.800 30.200 ;
        RECT 50.200 28.000 50.600 30.200 ;
        RECT 54.200 27.900 54.600 30.200 ;
        RECT 56.900 28.900 57.400 30.200 ;
        RECT 58.600 28.900 59.000 30.200 ;
        RECT 61.400 28.000 61.800 30.200 ;
        RECT 63.000 27.900 63.400 30.200 ;
        RECT 64.600 27.900 65.000 30.200 ;
        RECT 66.200 27.900 66.600 30.200 ;
        RECT 67.800 27.900 68.200 30.200 ;
        RECT 69.400 27.900 69.800 30.200 ;
        RECT 70.200 27.900 70.600 30.200 ;
        RECT 71.800 27.900 72.200 30.200 ;
        RECT 73.400 27.900 73.800 30.200 ;
        RECT 75.000 27.900 75.400 30.200 ;
        RECT 76.600 27.900 77.000 30.200 ;
        RECT 78.300 29.900 78.700 30.200 ;
        RECT 78.200 28.200 78.700 29.900 ;
        RECT 81.300 28.200 81.800 30.200 ;
        RECT 83.800 28.900 84.200 30.200 ;
        RECT 84.600 28.900 85.000 30.200 ;
        RECT 86.700 27.900 87.100 30.200 ;
        RECT 87.800 28.900 88.200 30.200 ;
        RECT 89.400 28.900 89.800 30.200 ;
        RECT 90.200 28.900 90.600 30.200 ;
        RECT 93.400 28.300 93.800 30.200 ;
        RECT 95.000 28.900 95.400 30.200 ;
        RECT 97.100 27.900 97.500 30.200 ;
        RECT 100.600 26.900 101.000 30.200 ;
        RECT 103.000 28.900 103.400 30.200 ;
        RECT 105.100 27.900 105.500 30.200 ;
        RECT 108.600 26.900 109.000 30.200 ;
        RECT 110.200 28.900 110.600 30.200 ;
        RECT 111.000 28.900 111.400 30.200 ;
        RECT 112.600 28.900 113.000 30.200 ;
        RECT 113.400 28.900 113.800 30.200 ;
        RECT 115.000 28.100 115.400 30.200 ;
        RECT 119.800 29.100 120.200 30.200 ;
        RECT 121.400 28.900 121.800 30.200 ;
        RECT 123.800 28.300 124.200 30.200 ;
        RECT 126.200 28.900 126.600 30.200 ;
        RECT 127.800 28.900 128.200 30.200 ;
        RECT 128.800 27.900 129.200 30.200 ;
        RECT 131.800 27.900 132.200 30.200 ;
        RECT 132.600 28.900 133.000 30.200 ;
        RECT 134.200 28.900 134.600 30.200 ;
        RECT 137.400 26.900 137.800 30.200 ;
        RECT 139.000 28.300 139.400 30.200 ;
        RECT 143.000 27.900 143.400 30.200 ;
        RECT 143.800 26.900 144.200 30.200 ;
        RECT 148.600 28.300 149.000 30.200 ;
        RECT 1.400 10.800 1.800 13.100 ;
        RECT 4.100 10.800 4.600 12.100 ;
        RECT 5.800 10.800 6.200 12.100 ;
        RECT 8.600 10.800 9.000 13.000 ;
        RECT 10.200 10.800 10.600 12.100 ;
        RECT 12.600 11.100 13.100 12.800 ;
        RECT 12.700 10.800 13.100 11.100 ;
        RECT 15.700 10.800 16.200 12.800 ;
        RECT 18.200 10.800 18.600 13.100 ;
        RECT 20.900 10.800 21.400 12.100 ;
        RECT 22.600 10.800 23.000 12.100 ;
        RECT 25.400 10.800 25.800 13.000 ;
        RECT 27.800 11.100 28.300 12.800 ;
        RECT 27.900 10.800 28.300 11.100 ;
        RECT 30.900 10.800 31.400 12.800 ;
        RECT 33.400 10.800 33.800 13.100 ;
        RECT 36.100 10.800 36.600 12.100 ;
        RECT 37.800 10.800 38.200 12.100 ;
        RECT 40.600 10.800 41.000 13.000 ;
        RECT 43.300 10.800 43.700 13.000 ;
        RECT 45.400 10.800 45.800 12.100 ;
        RECT 47.000 10.800 47.400 12.100 ;
        RECT 47.800 10.800 48.200 12.100 ;
        RECT 49.400 10.800 49.800 12.100 ;
        RECT 52.600 10.800 53.000 13.100 ;
        RECT 55.300 10.800 55.800 12.100 ;
        RECT 57.000 10.800 57.400 12.100 ;
        RECT 59.800 10.800 60.200 13.000 ;
        RECT 62.200 10.800 62.600 13.100 ;
        RECT 64.900 10.800 65.400 12.100 ;
        RECT 66.600 10.800 67.000 12.100 ;
        RECT 69.400 10.800 69.800 13.000 ;
        RECT 71.000 10.800 71.400 13.100 ;
        RECT 73.400 10.800 73.800 12.100 ;
        RECT 75.000 10.800 75.400 12.100 ;
        RECT 75.800 10.800 76.200 12.100 ;
        RECT 78.200 10.800 78.600 12.700 ;
        RECT 80.600 10.800 81.000 12.100 ;
        RECT 82.200 10.800 82.600 12.100 ;
        RECT 84.100 10.800 84.500 13.000 ;
        RECT 87.300 10.800 87.700 13.000 ;
        RECT 90.200 10.800 90.600 12.100 ;
        RECT 91.000 10.800 91.400 12.100 ;
        RECT 93.100 10.800 93.500 13.100 ;
        RECT 94.200 10.800 94.600 14.100 ;
        RECT 97.400 10.800 97.800 12.100 ;
        RECT 99.000 10.800 99.400 12.100 ;
        RECT 102.200 10.800 102.600 12.100 ;
        RECT 105.400 10.800 105.800 14.100 ;
        RECT 107.000 10.800 107.400 12.100 ;
        RECT 109.400 10.800 109.800 12.700 ;
        RECT 112.300 10.800 112.700 13.000 ;
        RECT 115.000 10.800 115.400 12.100 ;
        RECT 116.600 10.800 117.000 11.900 ;
        RECT 120.600 10.800 121.000 12.100 ;
        RECT 122.700 10.800 123.100 13.100 ;
        RECT 123.800 10.800 124.200 12.100 ;
        RECT 125.400 10.800 125.800 12.100 ;
        RECT 126.200 10.800 126.600 14.100 ;
        RECT 130.200 10.800 130.700 12.800 ;
        RECT 133.300 11.100 133.800 12.800 ;
        RECT 133.300 10.800 133.700 11.100 ;
        RECT 135.800 10.800 136.200 13.100 ;
        RECT 138.500 10.800 139.000 12.100 ;
        RECT 140.200 10.800 140.600 12.100 ;
        RECT 143.000 10.800 143.400 13.000 ;
        RECT 145.400 10.800 145.800 13.100 ;
        RECT 147.800 10.800 148.200 12.700 ;
        RECT 0.200 10.200 151.800 10.800 ;
        RECT 1.500 9.900 1.900 10.200 ;
        RECT 1.400 8.200 1.900 9.900 ;
        RECT 4.500 8.200 5.000 10.200 ;
        RECT 6.200 7.900 6.600 10.200 ;
        RECT 10.200 8.300 10.600 10.200 ;
        RECT 12.600 8.200 13.100 10.200 ;
        RECT 15.700 9.900 16.100 10.200 ;
        RECT 15.700 8.200 16.200 9.900 ;
        RECT 19.000 8.300 19.400 10.200 ;
        RECT 21.400 8.900 21.800 10.200 ;
        RECT 23.100 9.900 23.500 10.200 ;
        RECT 23.000 8.200 23.500 9.900 ;
        RECT 26.100 8.200 26.600 10.200 ;
        RECT 29.400 8.300 29.800 10.200 ;
        RECT 31.000 8.900 31.400 10.200 ;
        RECT 32.600 8.900 33.000 10.200 ;
        RECT 34.200 8.900 34.600 10.200 ;
        RECT 35.900 9.900 36.300 10.200 ;
        RECT 35.800 8.200 36.300 9.900 ;
        RECT 38.900 8.200 39.400 10.200 ;
        RECT 41.400 7.900 41.800 10.200 ;
        RECT 44.100 8.900 44.600 10.200 ;
        RECT 45.800 8.900 46.200 10.200 ;
        RECT 48.600 8.000 49.000 10.200 ;
        RECT 52.600 7.900 53.000 10.200 ;
        RECT 55.300 8.900 55.800 10.200 ;
        RECT 57.000 8.900 57.400 10.200 ;
        RECT 59.800 8.000 60.200 10.200 ;
        RECT 62.200 7.900 62.600 10.200 ;
        RECT 64.600 8.000 65.000 10.200 ;
        RECT 67.400 8.900 67.800 10.200 ;
        RECT 69.000 8.900 69.500 10.200 ;
        RECT 71.800 7.900 72.200 10.200 ;
        RECT 74.200 7.900 74.600 10.200 ;
        RECT 76.600 8.000 77.000 10.200 ;
        RECT 79.400 8.900 79.800 10.200 ;
        RECT 81.000 8.900 81.500 10.200 ;
        RECT 83.800 7.900 84.200 10.200 ;
        RECT 86.200 7.900 86.600 10.200 ;
        RECT 88.900 8.900 89.400 10.200 ;
        RECT 90.600 8.900 91.000 10.200 ;
        RECT 93.400 8.000 93.800 10.200 ;
        RECT 95.800 7.900 96.200 10.200 ;
        RECT 99.800 7.900 100.200 10.200 ;
        RECT 102.500 8.900 103.000 10.200 ;
        RECT 104.200 8.900 104.600 10.200 ;
        RECT 107.000 8.000 107.400 10.200 ;
        RECT 109.400 7.900 109.800 10.200 ;
        RECT 111.800 7.900 112.200 10.200 ;
        RECT 114.500 8.900 115.000 10.200 ;
        RECT 116.200 8.900 116.600 10.200 ;
        RECT 119.000 8.000 119.400 10.200 ;
        RECT 121.400 7.900 121.800 10.200 ;
        RECT 123.800 7.900 124.200 10.200 ;
        RECT 126.500 8.900 127.000 10.200 ;
        RECT 128.200 8.900 128.600 10.200 ;
        RECT 131.000 8.000 131.400 10.200 ;
        RECT 133.400 7.900 133.800 10.200 ;
        RECT 135.800 7.900 136.200 10.200 ;
        RECT 138.500 8.900 139.000 10.200 ;
        RECT 140.200 8.900 140.600 10.200 ;
        RECT 143.000 8.000 143.400 10.200 ;
        RECT 145.400 7.900 145.800 10.200 ;
        RECT 148.600 7.900 149.000 10.200 ;
      LAYER via1 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 100.900 130.300 101.300 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 100.900 110.300 101.300 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 100.900 90.300 101.300 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 100.900 70.300 101.300 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 100.900 50.300 101.300 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 100.900 30.300 101.300 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 100.900 10.300 101.300 10.700 ;
      LAYER metal2 ;
        RECT 100.000 130.300 101.600 130.700 ;
        RECT 100.000 110.300 101.600 110.700 ;
        RECT 100.000 90.300 101.600 90.700 ;
        RECT 100.000 70.300 101.600 70.700 ;
        RECT 100.000 50.300 101.600 50.700 ;
        RECT 100.000 30.300 101.600 30.700 ;
        RECT 100.000 10.300 101.600 10.700 ;
      LAYER via2 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 100.900 130.300 101.300 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 100.900 110.300 101.300 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 100.900 90.300 101.300 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 100.900 70.300 101.300 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 100.900 50.300 101.300 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 100.900 30.300 101.300 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 100.900 10.300 101.300 10.700 ;
      LAYER metal3 ;
        RECT 100.000 130.300 101.600 130.700 ;
        RECT 100.000 110.300 101.600 110.700 ;
        RECT 100.000 90.300 101.600 90.700 ;
        RECT 100.000 70.300 101.600 70.700 ;
        RECT 100.000 50.300 101.600 50.700 ;
        RECT 100.000 30.300 101.600 30.700 ;
        RECT 100.000 10.300 101.600 10.700 ;
      LAYER via3 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 101.000 130.300 101.400 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 101.000 110.300 101.400 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 101.000 90.300 101.400 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 101.000 70.300 101.400 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 101.000 50.300 101.400 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 101.000 30.300 101.400 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 101.000 10.300 101.400 10.700 ;
      LAYER metal4 ;
        RECT 100.000 130.300 101.600 130.700 ;
        RECT 100.000 110.300 101.600 110.700 ;
        RECT 100.000 90.300 101.600 90.700 ;
        RECT 100.000 70.300 101.600 70.700 ;
        RECT 100.000 50.300 101.600 50.700 ;
        RECT 100.000 30.300 101.600 30.700 ;
        RECT 100.000 10.300 101.600 10.700 ;
      LAYER via4 ;
        RECT 100.200 130.300 100.600 130.700 ;
        RECT 100.900 130.300 101.300 130.700 ;
        RECT 100.200 110.300 100.600 110.700 ;
        RECT 100.900 110.300 101.300 110.700 ;
        RECT 100.200 90.300 100.600 90.700 ;
        RECT 100.900 90.300 101.300 90.700 ;
        RECT 100.200 70.300 100.600 70.700 ;
        RECT 100.900 70.300 101.300 70.700 ;
        RECT 100.200 50.300 100.600 50.700 ;
        RECT 100.900 50.300 101.300 50.700 ;
        RECT 100.200 30.300 100.600 30.700 ;
        RECT 100.900 30.300 101.300 30.700 ;
        RECT 100.200 10.300 100.600 10.700 ;
        RECT 100.900 10.300 101.300 10.700 ;
      LAYER metal5 ;
        RECT 100.000 130.200 101.600 130.700 ;
        RECT 100.000 110.200 101.600 110.700 ;
        RECT 100.000 90.200 101.600 90.700 ;
        RECT 100.000 70.200 101.600 70.700 ;
        RECT 100.000 50.200 101.600 50.700 ;
        RECT 100.000 30.200 101.600 30.700 ;
        RECT 100.000 10.200 101.600 10.700 ;
      LAYER via5 ;
        RECT 101.000 130.200 101.500 130.700 ;
        RECT 101.000 110.200 101.500 110.700 ;
        RECT 101.000 90.200 101.500 90.700 ;
        RECT 101.000 70.200 101.500 70.700 ;
        RECT 101.000 50.200 101.500 50.700 ;
        RECT 101.000 30.200 101.500 30.700 ;
        RECT 101.000 10.200 101.500 10.700 ;
      LAYER metal6 ;
        RECT 100.000 -3.000 101.600 133.000 ;
    END
  END gnd
  PIN A[0]
    PORT
      LAYER metal1 ;
        RECT 45.200 126.900 45.600 127.000 ;
        RECT 45.200 126.600 45.700 126.900 ;
        RECT 45.400 126.200 45.700 126.600 ;
        RECT 45.400 125.800 45.800 126.200 ;
        RECT 47.000 125.400 47.400 126.200 ;
      LAYER via1 ;
        RECT 47.000 125.800 47.400 126.200 ;
      LAYER metal2 ;
        RECT 45.400 132.800 45.800 133.200 ;
        RECT 45.400 126.200 45.700 132.800 ;
        RECT 45.400 125.800 45.800 126.200 ;
        RECT 46.200 126.100 46.600 126.200 ;
        RECT 47.000 126.100 47.400 126.200 ;
        RECT 46.200 125.800 47.400 126.100 ;
      LAYER metal3 ;
        RECT 45.400 126.100 45.800 126.200 ;
        RECT 46.200 126.100 46.600 126.200 ;
        RECT 45.400 125.800 46.600 126.100 ;
    END
  END A[0]
  PIN A[1]
    PORT
      LAYER metal1 ;
        RECT 21.400 127.800 21.800 128.600 ;
        RECT 23.800 126.800 24.600 127.200 ;
      LAYER metal2 ;
        RECT 21.400 132.800 21.800 133.200 ;
        RECT 21.400 128.200 21.700 132.800 ;
        RECT 21.400 127.800 21.800 128.200 ;
        RECT 23.800 127.800 24.200 128.200 ;
        RECT 23.800 127.200 24.100 127.800 ;
        RECT 23.800 126.800 24.200 127.200 ;
      LAYER metal3 ;
        RECT 21.400 128.100 21.800 128.200 ;
        RECT 23.800 128.100 24.200 128.200 ;
        RECT 21.400 127.800 24.200 128.100 ;
    END
  END A[1]
  PIN A[2]
    PORT
      LAYER metal1 ;
        RECT 4.000 126.900 4.400 127.000 ;
        RECT 3.900 126.600 4.400 126.900 ;
        RECT 3.900 126.200 4.200 126.600 ;
        RECT 0.600 125.400 1.000 126.200 ;
        RECT 3.800 125.800 4.200 126.200 ;
      LAYER via1 ;
        RECT 0.600 125.800 1.000 126.200 ;
      LAYER metal2 ;
        RECT 0.600 125.800 1.000 126.200 ;
        RECT 3.800 125.800 4.200 126.200 ;
        RECT 0.600 125.200 0.900 125.800 ;
        RECT 3.800 125.200 4.100 125.800 ;
        RECT 0.600 124.800 1.000 125.200 ;
        RECT 3.800 124.800 4.200 125.200 ;
      LAYER metal3 ;
        RECT -2.600 125.100 -2.200 125.200 ;
        RECT 0.600 125.100 1.000 125.200 ;
        RECT 3.800 125.100 4.200 125.200 ;
        RECT -2.600 124.800 4.200 125.100 ;
    END
  END A[2]
  PIN A[3]
    PORT
      LAYER metal1 ;
        RECT 4.600 107.800 5.000 108.600 ;
        RECT 2.200 105.400 2.600 106.200 ;
      LAYER via1 ;
        RECT 2.200 105.800 2.600 106.200 ;
      LAYER metal2 ;
        RECT 4.600 107.800 5.000 108.200 ;
        RECT 2.200 105.800 2.600 106.200 ;
        RECT 2.200 105.200 2.500 105.800 ;
        RECT 4.600 105.200 4.900 107.800 ;
        RECT 2.200 104.800 2.600 105.200 ;
        RECT 4.600 104.800 5.000 105.200 ;
      LAYER metal3 ;
        RECT -2.600 105.100 -2.200 105.200 ;
        RECT 2.200 105.100 2.600 105.200 ;
        RECT 4.600 105.100 5.000 105.200 ;
        RECT -2.600 104.800 5.000 105.100 ;
    END
  END A[3]
  PIN A[4]
    PORT
      LAYER metal1 ;
        RECT 2.200 115.800 2.600 116.600 ;
        RECT 2.200 114.100 2.600 114.200 ;
        RECT 3.000 114.100 3.800 114.200 ;
        RECT 2.200 113.800 3.800 114.100 ;
      LAYER metal2 ;
        RECT 2.200 116.800 2.600 117.200 ;
        RECT 2.200 116.200 2.500 116.800 ;
        RECT 2.200 115.800 2.600 116.200 ;
        RECT 2.200 114.200 2.500 115.800 ;
        RECT 2.200 113.800 2.600 114.200 ;
      LAYER metal3 ;
        RECT -2.600 117.100 -2.200 117.200 ;
        RECT 2.200 117.100 2.600 117.200 ;
        RECT -2.600 116.800 2.600 117.100 ;
    END
  END A[4]
  PIN A[5]
    PORT
      LAYER metal1 ;
        RECT 2.200 73.800 2.600 74.200 ;
        RECT 2.200 73.200 2.500 73.800 ;
        RECT 2.200 72.400 2.600 73.200 ;
        RECT 2.200 65.400 2.600 66.200 ;
      LAYER via1 ;
        RECT 2.200 65.800 2.600 66.200 ;
      LAYER metal2 ;
        RECT 2.200 73.800 2.600 74.200 ;
        RECT 2.200 73.200 2.500 73.800 ;
        RECT 2.200 72.800 2.600 73.200 ;
        RECT 1.400 66.100 1.800 66.200 ;
        RECT 2.200 66.100 2.600 66.200 ;
        RECT 1.400 65.800 2.600 66.100 ;
      LAYER metal3 ;
        RECT 0.600 73.100 1.000 73.200 ;
        RECT 2.200 73.100 2.600 73.200 ;
        RECT 0.600 72.800 2.600 73.100 ;
        RECT -2.600 66.100 -2.200 66.200 ;
        RECT 0.600 66.100 1.000 66.200 ;
        RECT 1.400 66.100 1.800 66.200 ;
        RECT -2.600 65.800 1.800 66.100 ;
      LAYER via3 ;
        RECT 0.600 65.800 1.000 66.200 ;
      LAYER metal4 ;
        RECT 0.600 72.800 1.000 73.200 ;
        RECT 0.600 66.200 0.900 72.800 ;
        RECT 0.600 65.800 1.000 66.200 ;
    END
  END A[5]
  PIN A[6]
    PORT
      LAYER metal1 ;
        RECT 2.200 47.100 2.600 47.200 ;
        RECT 3.000 47.100 3.800 47.200 ;
        RECT 2.200 46.800 3.800 47.100 ;
        RECT 2.200 44.400 2.600 45.200 ;
      LAYER via1 ;
        RECT 2.200 44.800 2.600 45.200 ;
      LAYER metal2 ;
        RECT 2.200 46.800 2.600 47.200 ;
        RECT 2.200 45.200 2.500 46.800 ;
        RECT 2.200 44.800 2.600 45.200 ;
      LAYER metal3 ;
        RECT -2.600 45.100 -2.200 45.200 ;
        RECT 2.200 45.100 2.600 45.200 ;
        RECT -2.600 44.800 2.600 45.100 ;
    END
  END A[6]
  PIN A[7]
    PORT
      LAYER metal1 ;
        RECT 3.000 66.800 3.800 67.200 ;
      LAYER metal2 ;
        RECT 3.000 68.800 3.400 69.200 ;
        RECT 3.000 67.200 3.300 68.800 ;
        RECT 3.000 66.800 3.400 67.200 ;
      LAYER metal3 ;
        RECT 3.000 69.100 3.400 69.200 ;
        RECT -2.600 68.800 3.400 69.100 ;
        RECT -2.600 68.200 -2.300 68.800 ;
        RECT -2.600 67.800 -2.200 68.200 ;
    END
  END A[7]
  PIN B[0]
    PORT
      LAYER metal1 ;
        RECT 48.600 127.800 49.000 128.600 ;
        RECT 46.200 127.100 46.600 127.200 ;
        RECT 47.000 127.100 47.400 127.200 ;
        RECT 46.200 126.800 47.400 127.100 ;
        RECT 46.200 126.400 46.600 126.800 ;
      LAYER via1 ;
        RECT 47.000 126.800 47.400 127.200 ;
      LAYER metal2 ;
        RECT 47.800 133.100 48.200 133.200 ;
        RECT 47.000 132.800 48.200 133.100 ;
        RECT 47.000 128.200 47.300 132.800 ;
        RECT 47.000 127.800 47.400 128.200 ;
        RECT 47.800 128.100 48.200 128.200 ;
        RECT 48.600 128.100 49.000 128.200 ;
        RECT 47.800 127.800 49.000 128.100 ;
        RECT 47.000 127.200 47.300 127.800 ;
        RECT 47.000 126.800 47.400 127.200 ;
      LAYER metal3 ;
        RECT 47.000 128.100 47.400 128.200 ;
        RECT 47.800 128.100 48.200 128.200 ;
        RECT 47.000 127.800 48.200 128.100 ;
    END
  END B[0]
  PIN B[1]
    PORT
      LAYER metal1 ;
        RECT 23.000 127.800 23.400 128.600 ;
        RECT 28.200 127.100 29.000 127.200 ;
        RECT 27.900 127.000 29.000 127.100 ;
        RECT 26.800 126.800 29.000 127.000 ;
        RECT 26.800 126.700 28.200 126.800 ;
        RECT 26.800 126.600 27.200 126.700 ;
      LAYER via1 ;
        RECT 28.600 126.800 29.000 127.200 ;
      LAYER metal2 ;
        RECT 23.800 132.800 24.200 133.200 ;
        RECT 23.800 130.200 24.100 132.800 ;
        RECT 23.800 130.100 24.200 130.200 ;
        RECT 23.000 129.800 24.200 130.100 ;
        RECT 28.600 129.800 29.000 130.200 ;
        RECT 23.000 128.200 23.300 129.800 ;
        RECT 23.000 127.800 23.400 128.200 ;
        RECT 28.600 127.200 28.900 129.800 ;
        RECT 28.600 126.800 29.000 127.200 ;
      LAYER via2 ;
        RECT 23.800 129.800 24.200 130.200 ;
      LAYER metal3 ;
        RECT 23.800 130.100 24.200 130.200 ;
        RECT 28.600 130.100 29.000 130.200 ;
        RECT 23.800 129.800 29.000 130.100 ;
    END
  END B[1]
  PIN B[2]
    PORT
      LAYER metal1 ;
        RECT 2.200 127.800 2.600 128.600 ;
        RECT 2.200 127.100 2.500 127.800 ;
        RECT 3.000 127.100 3.400 127.200 ;
        RECT 2.200 126.800 3.400 127.100 ;
        RECT 2.200 126.200 2.500 126.800 ;
        RECT 3.000 126.400 3.400 126.800 ;
        RECT 2.200 125.800 2.600 126.200 ;
      LAYER metal2 ;
        RECT 2.200 126.800 2.600 127.200 ;
        RECT 2.200 126.200 2.500 126.800 ;
        RECT 2.200 125.800 2.600 126.200 ;
      LAYER metal3 ;
        RECT -2.600 127.100 -2.200 127.200 ;
        RECT 2.200 127.100 2.600 127.200 ;
        RECT -2.600 126.800 2.600 127.100 ;
    END
  END B[2]
  PIN B[3]
    PORT
      LAYER metal1 ;
        RECT 0.600 107.800 1.000 108.600 ;
        RECT 2.200 108.100 2.600 108.200 ;
        RECT 3.000 108.100 3.400 108.600 ;
        RECT 2.200 107.800 3.400 108.100 ;
      LAYER metal2 ;
        RECT 0.600 107.800 1.000 108.200 ;
        RECT 2.200 107.800 2.600 108.200 ;
        RECT 0.600 107.200 0.900 107.800 ;
        RECT 2.200 107.200 2.500 107.800 ;
        RECT 0.600 106.800 1.000 107.200 ;
        RECT 2.200 106.800 2.600 107.200 ;
      LAYER metal3 ;
        RECT -2.600 107.100 -2.200 107.200 ;
        RECT 0.600 107.100 1.000 107.200 ;
        RECT 2.200 107.100 2.600 107.200 ;
        RECT -2.600 106.800 2.600 107.100 ;
    END
  END B[3]
  PIN B[4]
    PORT
      LAYER metal1 ;
        RECT 6.000 114.300 6.400 114.400 ;
        RECT 6.000 114.200 7.400 114.300 ;
        RECT 0.600 113.400 1.000 114.200 ;
        RECT 6.000 114.000 8.200 114.200 ;
        RECT 7.100 113.900 8.200 114.000 ;
        RECT 7.400 113.800 8.200 113.900 ;
      LAYER via1 ;
        RECT 0.600 113.800 1.000 114.200 ;
        RECT 7.800 113.800 8.200 114.200 ;
      LAYER metal2 ;
        RECT 0.600 114.800 1.000 115.200 ;
        RECT 7.800 114.800 8.200 115.200 ;
        RECT 0.600 114.200 0.900 114.800 ;
        RECT 7.800 114.200 8.100 114.800 ;
        RECT 0.600 113.800 1.000 114.200 ;
        RECT 7.800 113.800 8.200 114.200 ;
      LAYER metal3 ;
        RECT -2.600 115.100 -2.200 115.200 ;
        RECT 0.600 115.100 1.000 115.200 ;
        RECT 7.800 115.100 8.200 115.200 ;
        RECT -2.600 114.800 8.200 115.100 ;
    END
  END B[4]
  PIN B[5]
    PORT
      LAYER metal1 ;
        RECT 0.600 72.400 1.000 73.200 ;
        RECT 0.600 67.800 1.000 68.600 ;
      LAYER via1 ;
        RECT 0.600 72.800 1.000 73.200 ;
      LAYER metal2 ;
        RECT 0.600 77.800 1.000 78.200 ;
        RECT 0.600 73.200 0.900 77.800 ;
        RECT 0.600 72.800 1.000 73.200 ;
        RECT 0.600 68.200 0.900 72.800 ;
        RECT 0.600 67.800 1.000 68.200 ;
      LAYER metal3 ;
        RECT -2.600 78.100 -2.200 78.200 ;
        RECT 0.600 78.100 1.000 78.200 ;
        RECT -2.600 77.800 1.000 78.100 ;
    END
  END B[5]
  PIN B[6]
    PORT
      LAYER metal1 ;
        RECT 0.600 46.800 1.000 47.600 ;
        RECT 4.500 47.400 4.900 47.800 ;
        RECT 5.800 47.700 6.600 47.800 ;
        RECT 5.800 47.400 6.800 47.700 ;
        RECT 4.500 47.200 4.800 47.400 ;
        RECT 4.400 46.800 4.800 47.200 ;
        RECT 6.500 47.200 6.800 47.400 ;
        RECT 6.500 46.900 8.200 47.200 ;
        RECT 7.400 46.800 8.200 46.900 ;
      LAYER via1 ;
        RECT 6.200 47.400 6.600 47.800 ;
      LAYER metal2 ;
        RECT 0.600 47.800 1.000 48.200 ;
        RECT 4.600 47.800 5.000 48.200 ;
        RECT 0.600 47.200 0.900 47.800 ;
        RECT 4.500 47.500 6.600 47.800 ;
        RECT 4.500 47.400 4.900 47.500 ;
        RECT 6.200 47.400 6.600 47.500 ;
        RECT 0.600 46.800 1.000 47.200 ;
      LAYER metal3 ;
        RECT 0.600 48.100 1.000 48.200 ;
        RECT 4.600 48.100 5.000 48.200 ;
        RECT 0.600 47.800 5.000 48.100 ;
        RECT -2.600 47.100 -2.200 47.200 ;
        RECT 0.600 47.100 1.000 47.200 ;
        RECT -2.600 46.800 1.000 47.100 ;
    END
  END B[6]
  PIN B[7]
    PORT
      LAYER metal1 ;
        RECT 4.500 67.400 4.900 67.800 ;
        RECT 5.800 67.700 6.600 67.800 ;
        RECT 5.800 67.400 6.800 67.700 ;
        RECT 4.500 67.200 4.800 67.400 ;
        RECT 4.400 66.800 4.800 67.200 ;
        RECT 6.500 67.200 6.800 67.400 ;
        RECT 6.500 66.900 8.200 67.200 ;
        RECT 7.400 66.800 8.200 66.900 ;
      LAYER via1 ;
        RECT 6.200 67.400 6.600 67.800 ;
      LAYER metal2 ;
        RECT 4.600 67.800 5.000 68.200 ;
        RECT 4.500 67.500 6.600 67.800 ;
        RECT 4.500 67.400 4.900 67.500 ;
        RECT 6.200 67.400 6.600 67.500 ;
      LAYER metal3 ;
        RECT -2.600 70.100 -2.200 70.200 ;
        RECT 1.400 70.100 1.800 70.200 ;
        RECT -2.600 69.800 1.800 70.100 ;
        RECT 1.400 68.100 1.800 68.200 ;
        RECT 4.600 68.100 5.000 68.200 ;
        RECT 1.400 67.800 5.000 68.100 ;
      LAYER via3 ;
        RECT 1.400 69.800 1.800 70.200 ;
      LAYER metal4 ;
        RECT 1.400 69.800 1.800 70.200 ;
        RECT 1.400 68.200 1.700 69.800 ;
        RECT 1.400 67.800 1.800 68.200 ;
    END
  END B[7]
  PIN C[0]
    PORT
      LAYER metal1 ;
        RECT 32.600 7.800 33.000 8.600 ;
        RECT 29.800 7.200 30.200 7.400 ;
        RECT 29.800 6.900 30.600 7.200 ;
        RECT 30.200 6.800 30.600 6.900 ;
        RECT 35.000 7.100 35.800 7.200 ;
        RECT 35.000 7.000 36.100 7.100 ;
        RECT 35.000 6.800 37.200 7.000 ;
        RECT 35.800 6.700 37.200 6.800 ;
        RECT 36.800 6.600 37.200 6.700 ;
      LAYER metal2 ;
        RECT 30.200 7.800 30.600 8.200 ;
        RECT 32.600 8.100 33.000 8.200 ;
        RECT 33.400 8.100 33.800 8.200 ;
        RECT 32.600 7.800 33.800 8.100 ;
        RECT 35.000 7.800 35.400 8.200 ;
        RECT 30.200 7.200 30.500 7.800 ;
        RECT 35.000 7.200 35.300 7.800 ;
        RECT 30.200 6.800 30.600 7.200 ;
        RECT 35.000 6.800 35.400 7.200 ;
        RECT 35.000 -1.900 35.300 6.800 ;
        RECT 35.800 -1.900 36.200 -1.800 ;
        RECT 35.000 -2.200 36.200 -1.900 ;
      LAYER via2 ;
        RECT 33.400 7.800 33.800 8.200 ;
      LAYER metal3 ;
        RECT 30.200 8.100 30.600 8.200 ;
        RECT 33.400 8.100 33.800 8.200 ;
        RECT 35.000 8.100 35.400 8.200 ;
        RECT 30.200 7.800 35.400 8.100 ;
    END
  END C[0]
  PIN C[1]
    PORT
      LAYER metal1 ;
        RECT 21.400 7.800 21.800 8.600 ;
        RECT 21.400 7.100 21.700 7.800 ;
        RECT 23.800 7.700 24.600 7.800 ;
        RECT 23.600 7.400 24.600 7.700 ;
        RECT 25.500 7.400 25.900 7.800 ;
        RECT 23.600 7.200 23.900 7.400 ;
        RECT 22.200 7.100 23.900 7.200 ;
        RECT 21.400 6.900 23.900 7.100 ;
        RECT 25.600 7.200 25.900 7.400 ;
        RECT 21.400 6.800 23.000 6.900 ;
        RECT 25.600 6.800 26.000 7.200 ;
      LAYER via1 ;
        RECT 23.800 7.400 24.200 7.800 ;
        RECT 22.200 6.800 22.600 7.200 ;
      LAYER metal2 ;
        RECT 23.800 7.500 25.900 7.800 ;
        RECT 23.800 7.400 24.200 7.500 ;
        RECT 25.500 7.400 25.900 7.500 ;
        RECT 22.200 6.800 22.600 7.200 ;
        RECT 22.200 -1.900 22.500 6.800 ;
        RECT 23.800 -1.900 24.200 -1.800 ;
        RECT 22.200 -2.200 24.200 -1.900 ;
    END
  END C[1]
  PIN C[2]
    PORT
      LAYER metal1 ;
        RECT 11.800 14.100 12.600 14.200 ;
        RECT 11.800 13.800 13.500 14.100 ;
        RECT 13.200 13.600 13.500 13.800 ;
        RECT 15.200 13.800 15.600 14.200 ;
        RECT 15.200 13.600 15.500 13.800 ;
        RECT 13.200 13.300 14.200 13.600 ;
        RECT 13.400 13.200 14.200 13.300 ;
        RECT 15.100 13.200 15.500 13.600 ;
        RECT 10.200 12.400 10.600 13.200 ;
      LAYER via1 ;
        RECT 10.200 12.800 10.600 13.200 ;
      LAYER metal2 ;
        RECT 13.400 13.500 13.800 13.600 ;
        RECT 15.100 13.500 15.500 13.600 ;
        RECT 13.400 13.200 15.500 13.500 ;
        RECT 10.200 13.100 10.600 13.200 ;
        RECT 11.000 13.100 11.400 13.200 ;
        RECT 10.200 12.800 11.400 13.100 ;
        RECT 13.400 12.800 13.800 13.200 ;
      LAYER via2 ;
        RECT 11.000 12.800 11.400 13.200 ;
      LAYER metal3 ;
        RECT -2.600 13.100 -2.200 13.200 ;
        RECT 11.000 13.100 11.400 13.200 ;
        RECT 13.400 13.100 13.800 13.200 ;
        RECT -2.600 12.800 13.800 13.100 ;
    END
  END C[2]
  PIN C[3]
    PORT
      LAYER metal1 ;
        RECT 6.200 74.100 7.000 74.200 ;
        RECT 5.400 73.800 7.900 74.100 ;
        RECT 5.400 73.200 5.700 73.800 ;
        RECT 7.600 73.600 7.900 73.800 ;
        RECT 9.600 73.800 10.000 74.200 ;
        RECT 9.600 73.600 9.900 73.800 ;
        RECT 7.600 73.300 8.600 73.600 ;
        RECT 7.800 73.200 8.600 73.300 ;
        RECT 9.500 73.200 9.900 73.600 ;
        RECT 5.400 72.800 5.800 73.200 ;
        RECT 11.800 72.400 12.200 73.200 ;
      LAYER via1 ;
        RECT 11.800 72.800 12.200 73.200 ;
      LAYER metal2 ;
        RECT 5.400 73.800 5.800 74.200 ;
        RECT 5.400 73.200 5.700 73.800 ;
        RECT 7.800 73.500 8.200 73.600 ;
        RECT 9.500 73.500 9.900 73.600 ;
        RECT 7.800 73.200 9.900 73.500 ;
        RECT 5.400 72.800 5.800 73.200 ;
        RECT 9.400 72.800 9.800 73.200 ;
        RECT 11.000 73.100 11.400 73.200 ;
        RECT 11.800 73.100 12.200 73.200 ;
        RECT 11.000 72.800 12.200 73.100 ;
      LAYER metal3 ;
        RECT -2.600 74.100 -2.200 74.200 ;
        RECT 5.400 74.100 5.800 74.200 ;
        RECT -2.600 73.800 5.800 74.100 ;
        RECT 9.400 73.100 9.800 73.200 ;
        RECT 11.000 73.100 11.400 73.200 ;
        RECT 9.400 72.800 11.400 73.100 ;
    END
  END C[3]
  PIN C[4]
    PORT
      LAYER metal1 ;
        RECT 0.600 92.400 1.000 93.200 ;
      LAYER via1 ;
        RECT 0.600 92.800 1.000 93.200 ;
      LAYER metal2 ;
        RECT 0.600 94.800 1.000 95.200 ;
        RECT 0.600 93.200 0.900 94.800 ;
        RECT 0.600 92.800 1.000 93.200 ;
      LAYER metal3 ;
        RECT -2.600 95.100 -2.200 95.200 ;
        RECT 0.600 95.100 1.000 95.200 ;
        RECT -2.600 94.800 1.000 95.100 ;
    END
  END C[4]
  PIN C[5]
    PORT
      LAYER metal1 ;
        RECT 0.600 87.800 1.000 88.600 ;
      LAYER metal2 ;
        RECT 0.600 87.800 1.000 88.200 ;
        RECT 0.600 87.200 0.900 87.800 ;
        RECT 0.600 86.800 1.000 87.200 ;
      LAYER metal3 ;
        RECT -2.600 87.100 -2.200 87.200 ;
        RECT 0.600 87.100 1.000 87.200 ;
        RECT -2.600 86.800 1.000 87.100 ;
    END
  END C[5]
  PIN C[6]
    PORT
      LAYER metal1 ;
        RECT 2.400 34.300 2.800 34.400 ;
        RECT 1.400 34.200 2.800 34.300 ;
        RECT 0.600 34.000 2.800 34.200 ;
        RECT 0.600 33.900 1.700 34.000 ;
        RECT 0.600 33.800 1.400 33.900 ;
        RECT 6.200 33.400 6.600 34.200 ;
      LAYER via1 ;
        RECT 6.200 33.800 6.600 34.200 ;
      LAYER metal2 ;
        RECT 0.600 35.800 1.000 36.200 ;
        RECT 6.200 35.800 6.600 36.200 ;
        RECT 0.600 34.200 0.900 35.800 ;
        RECT 6.200 34.200 6.500 35.800 ;
        RECT 0.600 33.800 1.000 34.200 ;
        RECT 6.200 33.800 6.600 34.200 ;
      LAYER metal3 ;
        RECT -2.600 36.100 -2.200 36.200 ;
        RECT 0.600 36.100 1.000 36.200 ;
        RECT 6.200 36.100 6.600 36.200 ;
        RECT -2.600 35.800 6.600 36.100 ;
    END
  END C[6]
  PIN C[7]
    PORT
      LAYER metal1 ;
        RECT 0.600 7.100 1.400 7.200 ;
        RECT 0.600 7.000 1.700 7.100 ;
        RECT 0.600 6.800 2.800 7.000 ;
        RECT 1.400 6.700 2.800 6.800 ;
        RECT 2.400 6.600 2.800 6.700 ;
      LAYER metal2 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 0.600 5.200 0.900 6.800 ;
        RECT 0.600 4.800 1.000 5.200 ;
      LAYER metal3 ;
        RECT -2.600 5.100 -2.200 5.200 ;
        RECT 0.600 5.100 1.000 5.200 ;
        RECT -2.600 4.800 1.000 5.100 ;
    END
  END C[7]
  PIN D[0]
    PORT
      LAYER metal1 ;
        RECT 34.200 7.800 34.600 8.600 ;
        RECT 39.400 6.800 40.200 7.200 ;
        RECT 41.700 6.200 42.100 6.300 ;
        RECT 43.000 6.200 43.400 6.300 ;
        RECT 41.700 5.900 44.200 6.200 ;
        RECT 43.800 5.800 44.200 5.900 ;
      LAYER via1 ;
        RECT 39.800 6.800 40.200 7.200 ;
        RECT 43.000 5.900 43.400 6.300 ;
      LAYER metal2 ;
        RECT 34.200 7.800 34.600 8.200 ;
        RECT 34.200 6.200 34.500 7.800 ;
        RECT 39.800 6.800 40.200 7.200 ;
        RECT 39.800 6.200 40.100 6.800 ;
        RECT 43.000 6.200 43.400 6.300 ;
        RECT 43.800 6.200 44.200 6.300 ;
        RECT 34.200 5.800 34.600 6.200 ;
        RECT 39.800 5.800 40.200 6.200 ;
        RECT 43.000 5.900 44.200 6.200 ;
        RECT 43.000 -1.800 43.300 5.900 ;
        RECT 43.000 -2.200 43.400 -1.800 ;
      LAYER via2 ;
        RECT 43.800 5.900 44.200 6.300 ;
      LAYER metal3 ;
        RECT 34.200 6.100 34.600 6.200 ;
        RECT 39.800 6.100 40.200 6.200 ;
        RECT 43.800 6.100 44.200 6.300 ;
        RECT 34.200 5.900 44.200 6.100 ;
        RECT 34.200 5.800 44.100 5.900 ;
    END
  END D[0]
  PIN D[1]
    PORT
      LAYER metal1 ;
        RECT 26.600 6.800 27.400 7.200 ;
        RECT 19.000 5.800 19.400 6.600 ;
        RECT 52.900 6.200 53.300 6.300 ;
        RECT 54.200 6.200 54.600 6.300 ;
        RECT 52.900 5.900 55.400 6.200 ;
        RECT 55.000 5.800 55.400 5.900 ;
      LAYER via1 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 54.200 5.900 54.600 6.300 ;
      LAYER metal2 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 55.000 6.800 55.400 7.200 ;
        RECT 27.000 6.200 27.300 6.800 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 19.800 6.100 20.200 6.200 ;
        RECT 19.000 5.800 20.200 6.100 ;
        RECT 27.000 5.800 27.400 6.200 ;
        RECT 54.200 5.900 54.600 6.300 ;
        RECT 55.000 6.200 55.300 6.800 ;
        RECT 54.200 -1.800 54.500 5.900 ;
        RECT 55.000 5.800 55.400 6.200 ;
        RECT 54.200 -2.200 54.600 -1.800 ;
      LAYER via2 ;
        RECT 19.800 5.800 20.200 6.200 ;
      LAYER metal3 ;
        RECT 27.000 7.100 27.400 7.200 ;
        RECT 55.000 7.100 55.400 7.200 ;
        RECT 27.000 6.800 55.400 7.100 ;
        RECT 19.800 6.100 20.200 6.200 ;
        RECT 27.000 6.100 27.400 6.200 ;
        RECT 19.800 5.800 27.400 6.100 ;
    END
  END D[1]
  PIN D[2]
    PORT
      LAYER metal1 ;
        RECT 20.600 15.100 21.000 15.200 ;
        RECT 18.500 14.800 21.000 15.100 ;
        RECT 18.500 14.700 18.900 14.800 ;
        RECT 19.800 14.700 20.200 14.800 ;
        RECT 16.200 13.800 17.000 14.200 ;
        RECT 10.200 5.800 10.600 6.600 ;
      LAYER via1 ;
        RECT 16.600 13.800 17.000 14.200 ;
      LAYER metal2 ;
        RECT 16.600 14.800 17.000 15.200 ;
        RECT 16.600 14.200 16.900 14.800 ;
        RECT 19.800 14.700 20.200 15.100 ;
        RECT 19.800 14.200 20.100 14.700 ;
        RECT 16.600 13.800 17.000 14.200 ;
        RECT 19.800 13.800 20.200 14.200 ;
        RECT 16.600 8.200 16.900 13.800 ;
        RECT 10.200 7.800 10.600 8.200 ;
        RECT 16.600 7.800 17.000 8.200 ;
        RECT 10.200 6.200 10.500 7.800 ;
        RECT 10.200 5.800 10.600 6.200 ;
        RECT 10.200 -1.800 10.500 5.800 ;
        RECT 10.200 -2.200 10.600 -1.800 ;
      LAYER metal3 ;
        RECT 16.600 15.100 17.000 15.200 ;
        RECT 16.600 14.800 20.100 15.100 ;
        RECT 19.800 14.200 20.100 14.800 ;
        RECT 19.800 13.800 20.200 14.200 ;
        RECT 10.200 8.100 10.600 8.200 ;
        RECT 16.600 8.100 17.000 8.200 ;
        RECT 10.200 7.800 17.000 8.100 ;
    END
  END D[2]
  PIN D[3]
    PORT
      LAYER metal1 ;
        RECT 14.200 74.400 14.600 75.200 ;
        RECT 23.000 75.100 23.400 75.200 ;
        RECT 20.900 74.800 23.400 75.100 ;
        RECT 20.900 74.700 21.300 74.800 ;
        RECT 22.200 74.700 22.600 74.800 ;
        RECT 10.600 74.100 11.400 74.200 ;
        RECT 11.800 74.100 12.200 74.200 ;
        RECT 10.600 73.800 12.200 74.100 ;
      LAYER via1 ;
        RECT 14.200 74.800 14.600 75.200 ;
        RECT 11.800 73.800 12.200 74.200 ;
      LAYER metal2 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 13.400 75.100 13.800 75.200 ;
        RECT 14.200 75.100 14.600 75.200 ;
        RECT 13.400 74.800 14.600 75.100 ;
        RECT 22.200 75.000 22.600 75.100 ;
        RECT 23.000 75.000 23.400 75.100 ;
        RECT 11.800 74.200 12.100 74.800 ;
        RECT 22.200 74.700 23.400 75.000 ;
        RECT 11.800 73.800 12.200 74.200 ;
      LAYER via2 ;
        RECT 23.000 74.700 23.400 75.100 ;
      LAYER metal3 ;
        RECT -2.600 76.100 -2.200 76.200 ;
        RECT -2.600 75.800 12.100 76.100 ;
        RECT 11.800 75.200 12.100 75.800 ;
        RECT 11.800 75.100 12.200 75.200 ;
        RECT 13.400 75.100 13.800 75.200 ;
        RECT 11.800 74.800 23.400 75.100 ;
        RECT 23.000 74.700 23.400 74.800 ;
    END
  END D[3]
  PIN D[4]
    PORT
      LAYER metal1 ;
        RECT 3.800 94.100 4.200 94.200 ;
        RECT 3.800 93.800 4.900 94.100 ;
        RECT 3.800 93.400 4.200 93.800 ;
        RECT 4.600 93.200 4.900 93.800 ;
        RECT 4.600 92.400 5.000 93.200 ;
        RECT 32.600 75.100 33.000 75.200 ;
        RECT 30.500 74.800 33.000 75.100 ;
        RECT 30.500 74.700 30.900 74.800 ;
        RECT 31.800 74.700 32.200 74.800 ;
      LAYER metal2 ;
        RECT 3.800 96.800 4.200 97.200 ;
        RECT 31.800 96.800 32.200 97.200 ;
        RECT 3.800 94.200 4.100 96.800 ;
        RECT 3.800 93.800 4.200 94.200 ;
        RECT 31.800 75.100 32.100 96.800 ;
        RECT 31.800 74.700 32.200 75.100 ;
      LAYER metal3 ;
        RECT -2.600 97.100 -2.200 97.200 ;
        RECT 3.800 97.100 4.200 97.200 ;
        RECT 31.800 97.100 32.200 97.200 ;
        RECT -2.600 96.800 32.200 97.100 ;
    END
  END D[4]
  PIN D[5]
    PORT
      LAYER metal1 ;
        RECT 2.200 86.800 2.600 87.600 ;
        RECT 5.400 86.800 5.900 87.200 ;
        RECT 2.200 86.200 2.500 86.800 ;
        RECT 5.600 86.400 6.000 86.800 ;
        RECT 39.300 86.200 39.700 86.300 ;
        RECT 40.600 86.200 41.000 86.300 ;
        RECT 2.200 85.800 2.600 86.200 ;
        RECT 39.300 85.900 41.800 86.200 ;
        RECT 41.400 85.800 41.800 85.900 ;
      LAYER via1 ;
        RECT 40.600 85.900 41.000 86.300 ;
      LAYER metal2 ;
        RECT 2.200 86.800 2.600 87.200 ;
        RECT 4.600 87.100 5.000 87.200 ;
        RECT 5.400 87.100 5.800 87.200 ;
        RECT 4.600 86.800 5.800 87.100 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 2.200 86.200 2.500 86.800 ;
        RECT 40.600 86.300 40.900 86.800 ;
        RECT 2.200 85.800 2.600 86.200 ;
        RECT 40.600 85.900 41.000 86.300 ;
      LAYER metal3 ;
        RECT 1.400 87.100 1.800 87.200 ;
        RECT 2.200 87.100 2.600 87.200 ;
        RECT 4.600 87.100 5.000 87.200 ;
        RECT 40.600 87.100 41.000 87.200 ;
        RECT 1.400 86.800 41.000 87.100 ;
        RECT -2.600 85.100 -2.200 85.200 ;
        RECT 1.400 85.100 1.800 85.200 ;
        RECT -2.600 84.800 1.800 85.100 ;
      LAYER via3 ;
        RECT 1.400 84.800 1.800 85.200 ;
      LAYER metal4 ;
        RECT 1.400 86.800 1.800 87.200 ;
        RECT 1.400 85.200 1.700 86.800 ;
        RECT 1.400 84.800 1.800 85.200 ;
    END
  END D[5]
  PIN D[6]
    PORT
      LAYER metal1 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 31.800 35.100 32.200 35.200 ;
        RECT 29.700 34.800 32.200 35.100 ;
        RECT 5.400 34.200 5.700 34.800 ;
        RECT 29.700 34.700 30.100 34.800 ;
        RECT 31.000 34.700 31.400 34.800 ;
        RECT 5.000 33.800 5.800 34.200 ;
        RECT 9.400 32.400 9.800 33.200 ;
      LAYER via1 ;
        RECT 9.400 32.800 9.800 33.200 ;
      LAYER metal2 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 5.400 34.200 5.700 34.800 ;
        RECT 31.000 34.700 31.400 35.100 ;
        RECT 31.000 34.200 31.300 34.700 ;
        RECT 5.400 33.800 5.800 34.200 ;
        RECT 9.400 33.800 9.800 34.200 ;
        RECT 31.000 33.800 31.400 34.200 ;
        RECT 9.400 33.200 9.700 33.800 ;
        RECT 9.400 32.800 9.800 33.200 ;
      LAYER metal3 ;
        RECT -2.600 34.100 -2.200 34.200 ;
        RECT 5.400 34.100 5.800 34.200 ;
        RECT 9.400 34.100 9.800 34.200 ;
        RECT 31.000 34.100 31.400 34.200 ;
        RECT -2.600 33.800 31.400 34.100 ;
    END
  END D[6]
  PIN D[7]
    PORT
      LAYER metal1 ;
        RECT 3.800 15.100 4.200 15.200 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 1.700 14.800 5.800 15.100 ;
        RECT 1.700 14.700 2.100 14.800 ;
        RECT 5.000 6.800 5.800 7.200 ;
      LAYER via1 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 5.400 6.800 5.800 7.200 ;
      LAYER metal2 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 5.400 7.200 5.700 14.800 ;
        RECT 5.400 6.800 5.800 7.200 ;
      LAYER metal3 ;
        RECT -2.600 15.100 -2.200 15.200 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT -2.600 14.800 5.800 15.100 ;
    END
  END D[7]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 37.700 54.100 38.600 54.500 ;
        RECT 38.200 53.800 38.600 54.100 ;
        RECT 33.400 46.900 33.800 47.200 ;
        RECT 73.400 46.900 73.800 47.200 ;
        RECT 32.900 46.500 33.800 46.900 ;
        RECT 72.900 46.500 73.800 46.900 ;
        RECT 0.600 26.900 1.000 27.200 ;
        RECT 69.400 27.100 69.800 27.200 ;
        RECT 70.200 27.100 70.600 27.200 ;
        RECT 69.400 26.900 70.600 27.100 ;
        RECT 0.600 26.500 1.500 26.900 ;
        RECT 68.900 26.800 71.100 26.900 ;
        RECT 68.900 26.500 69.800 26.800 ;
        RECT 70.200 26.500 71.100 26.800 ;
      LAYER via1 ;
        RECT 33.400 46.800 33.800 47.200 ;
        RECT 73.400 46.800 73.800 47.200 ;
        RECT 0.600 26.800 1.000 27.200 ;
        RECT 70.200 26.800 70.600 27.200 ;
      LAYER metal2 ;
        RECT 38.200 53.800 38.600 54.200 ;
        RECT 38.200 53.200 38.500 53.800 ;
        RECT 33.400 52.800 33.800 53.200 ;
        RECT 38.200 52.800 38.600 53.200 ;
        RECT 33.400 47.200 33.700 52.800 ;
        RECT 33.400 46.800 33.800 47.200 ;
        RECT 73.400 46.800 73.800 47.200 ;
        RECT 33.400 44.200 33.700 46.800 ;
        RECT 73.400 45.200 73.700 46.800 ;
        RECT 70.200 44.800 70.600 45.200 ;
        RECT 73.400 44.800 73.800 45.200 ;
        RECT 70.200 44.200 70.500 44.800 ;
        RECT 33.400 43.800 33.800 44.200 ;
        RECT 70.200 43.800 70.600 44.200 ;
        RECT 70.200 27.200 70.500 43.800 ;
        RECT 0.600 27.100 1.000 27.200 ;
        RECT 1.400 27.100 1.800 27.200 ;
        RECT 0.600 26.800 1.800 27.100 ;
        RECT 70.200 26.800 70.600 27.200 ;
      LAYER via2 ;
        RECT 1.400 26.800 1.800 27.200 ;
      LAYER metal3 ;
        RECT 33.400 53.100 33.800 53.200 ;
        RECT 38.200 53.100 38.600 53.200 ;
        RECT 33.400 52.800 38.600 53.100 ;
        RECT 70.200 45.100 70.600 45.200 ;
        RECT 73.400 45.100 73.800 45.200 ;
        RECT 70.200 44.800 73.800 45.100 ;
        RECT 0.600 44.100 1.000 44.200 ;
        RECT 33.400 44.100 33.800 44.200 ;
        RECT 70.200 44.100 70.600 44.200 ;
        RECT 0.600 43.800 70.600 44.100 ;
        RECT -2.600 27.100 -2.200 27.200 ;
        RECT 0.600 27.100 1.000 27.200 ;
        RECT 1.400 27.100 1.800 27.200 ;
        RECT -2.600 26.800 1.800 27.100 ;
      LAYER via3 ;
        RECT 0.600 26.800 1.000 27.200 ;
      LAYER metal4 ;
        RECT 0.600 43.800 1.000 44.200 ;
        RECT 0.600 27.200 0.900 43.800 ;
        RECT 0.600 26.800 1.000 27.200 ;
    END
  END clk
  PIN F[0]
    PORT
      LAYER metal1 ;
        RECT 61.400 6.200 61.800 9.900 ;
        RECT 61.400 5.100 61.700 6.200 ;
        RECT 61.400 1.100 61.800 5.100 ;
      LAYER via1 ;
        RECT 61.400 1.800 61.800 2.200 ;
      LAYER metal2 ;
        RECT 61.400 1.800 61.800 2.200 ;
        RECT 61.400 -1.900 61.700 1.800 ;
        RECT 62.200 -1.900 62.600 -1.800 ;
        RECT 61.400 -2.200 62.600 -1.900 ;
    END
  END F[0]
  PIN F[1]
    PORT
      LAYER metal1 ;
        RECT 73.400 6.200 73.800 9.900 ;
        RECT 73.400 5.100 73.700 6.200 ;
        RECT 73.400 1.100 73.800 5.100 ;
      LAYER via1 ;
        RECT 73.400 1.800 73.800 2.200 ;
      LAYER metal2 ;
        RECT 73.400 1.800 73.800 2.200 ;
        RECT 73.400 -1.900 73.700 1.800 ;
        RECT 74.200 -1.900 74.600 -1.800 ;
        RECT 73.400 -2.200 74.600 -1.900 ;
    END
  END F[1]
  PIN F[2]
    PORT
      LAYER metal1 ;
        RECT 96.600 6.200 97.000 9.900 ;
        RECT 96.700 5.100 97.000 6.200 ;
        RECT 96.600 1.100 97.000 5.100 ;
      LAYER via1 ;
        RECT 96.600 1.800 97.000 2.200 ;
      LAYER metal2 ;
        RECT 96.600 1.800 97.000 2.200 ;
        RECT 95.800 -1.900 96.200 -1.800 ;
        RECT 96.600 -1.900 96.900 1.800 ;
        RECT 95.800 -2.200 96.900 -1.900 ;
    END
  END F[2]
  PIN F[3]
    PORT
      LAYER metal1 ;
        RECT 110.200 6.200 110.600 9.900 ;
        RECT 110.300 5.100 110.600 6.200 ;
        RECT 110.200 1.100 110.600 5.100 ;
      LAYER via1 ;
        RECT 110.200 1.800 110.600 2.200 ;
      LAYER metal2 ;
        RECT 110.200 1.800 110.600 2.200 ;
        RECT 109.400 -1.900 109.800 -1.800 ;
        RECT 110.200 -1.900 110.500 1.800 ;
        RECT 109.400 -2.200 110.500 -1.900 ;
    END
  END F[3]
  PIN F[4]
    PORT
      LAYER metal1 ;
        RECT 122.200 6.200 122.600 9.900 ;
        RECT 122.300 5.100 122.600 6.200 ;
        RECT 122.200 1.100 122.600 5.100 ;
      LAYER via1 ;
        RECT 122.200 1.800 122.600 2.200 ;
      LAYER metal2 ;
        RECT 122.200 1.800 122.600 2.200 ;
        RECT 121.400 -1.900 121.800 -1.800 ;
        RECT 122.200 -1.900 122.500 1.800 ;
        RECT 121.400 -2.200 122.500 -1.900 ;
    END
  END F[4]
  PIN F[5]
    PORT
      LAYER metal1 ;
        RECT 134.200 6.200 134.600 9.900 ;
        RECT 134.300 5.100 134.600 6.200 ;
        RECT 134.200 1.100 134.600 5.100 ;
      LAYER via1 ;
        RECT 134.200 1.800 134.600 2.200 ;
      LAYER metal2 ;
        RECT 134.200 1.800 134.600 2.200 ;
        RECT 133.400 -1.900 133.800 -1.800 ;
        RECT 134.200 -1.900 134.500 1.800 ;
        RECT 133.400 -2.200 134.500 -1.900 ;
    END
  END F[5]
  PIN F[6]
    PORT
      LAYER metal1 ;
        RECT 146.200 15.900 146.600 19.900 ;
        RECT 146.300 14.800 146.600 15.900 ;
        RECT 146.200 11.100 146.600 14.800 ;
      LAYER via1 ;
        RECT 146.200 13.800 146.600 14.200 ;
      LAYER metal2 ;
        RECT 146.200 14.800 146.600 15.200 ;
        RECT 146.200 14.200 146.500 14.800 ;
        RECT 146.200 13.800 146.600 14.200 ;
      LAYER metal3 ;
        RECT 146.200 15.100 146.600 15.200 ;
        RECT 154.200 15.100 154.600 15.200 ;
        RECT 146.200 14.800 154.600 15.100 ;
    END
  END F[6]
  PIN F[7]
    PORT
      LAYER metal1 ;
        RECT 146.200 6.200 146.600 9.900 ;
        RECT 146.300 5.100 146.600 6.200 ;
        RECT 146.200 1.100 146.600 5.100 ;
      LAYER via1 ;
        RECT 146.200 1.800 146.600 2.200 ;
      LAYER metal2 ;
        RECT 146.200 1.800 146.600 2.200 ;
        RECT 145.400 -1.900 145.800 -1.800 ;
        RECT 146.200 -1.900 146.500 1.800 ;
        RECT 145.400 -2.200 146.500 -1.900 ;
    END
  END F[7]
  OBS
      LAYER metal1 ;
        RECT 1.400 128.900 1.800 129.900 ;
        RECT 0.600 128.100 1.000 128.200 ;
        RECT 1.400 128.100 1.700 128.900 ;
        RECT 0.600 127.800 1.700 128.100 ;
        RECT 3.000 127.900 3.400 129.900 ;
        RECT 5.100 128.400 5.500 129.900 ;
        RECT 7.000 128.900 7.400 129.900 ;
        RECT 5.100 127.900 5.800 128.400 ;
        RECT 1.400 127.200 1.700 127.800 ;
        RECT 3.100 127.800 3.400 127.900 ;
        RECT 3.100 127.600 4.000 127.800 ;
        RECT 3.100 127.500 5.200 127.600 ;
        RECT 3.700 127.300 5.200 127.500 ;
        RECT 4.800 127.200 5.200 127.300 ;
        RECT 1.400 126.800 1.800 127.200 ;
        RECT 1.400 125.100 1.700 126.800 ;
        RECT 4.800 125.500 5.100 127.200 ;
        RECT 5.500 126.200 5.800 127.900 ;
        RECT 6.200 127.800 6.600 128.600 ;
        RECT 7.100 127.200 7.400 128.900 ;
        RECT 8.700 128.200 9.100 128.600 ;
        RECT 7.800 128.100 8.200 128.200 ;
        RECT 8.600 128.100 9.000 128.200 ;
        RECT 7.800 127.800 9.000 128.100 ;
        RECT 9.400 127.900 9.800 129.900 ;
        RECT 5.400 126.100 5.800 126.200 ;
        RECT 6.200 126.800 6.600 127.200 ;
        RECT 7.000 127.100 7.400 127.200 ;
        RECT 8.600 127.100 9.000 127.200 ;
        RECT 7.000 126.800 9.000 127.100 ;
        RECT 6.200 126.100 6.500 126.800 ;
        RECT 5.400 125.800 6.500 126.100 ;
        RECT 3.900 125.200 5.100 125.500 ;
        RECT 0.900 124.700 1.800 125.100 ;
        RECT 0.900 121.100 1.300 124.700 ;
        RECT 3.900 123.100 4.200 125.200 ;
        RECT 5.500 125.100 5.800 125.800 ;
        RECT 7.100 125.100 7.400 126.800 ;
        RECT 9.500 126.200 9.800 127.900 ;
        RECT 11.800 127.900 12.200 129.900 ;
        RECT 14.000 128.100 14.800 129.900 ;
        RECT 11.800 127.600 13.000 127.900 ;
        RECT 12.600 127.500 13.000 127.600 ;
        RECT 13.300 127.400 13.700 127.800 ;
        RECT 13.300 127.200 13.600 127.400 ;
        RECT 10.200 126.400 10.600 127.200 ;
        RECT 11.800 126.800 12.600 127.200 ;
        RECT 13.200 126.800 13.600 127.200 ;
        RECT 14.000 127.100 14.300 128.100 ;
        RECT 16.600 127.900 17.000 129.900 ;
        RECT 17.400 127.900 17.800 129.900 ;
        RECT 18.200 128.000 18.600 129.900 ;
        RECT 19.800 128.000 20.200 129.900 ;
        RECT 18.200 127.900 20.200 128.000 ;
        RECT 14.600 127.400 15.400 127.800 ;
        RECT 15.700 127.600 17.000 127.900 ;
        RECT 15.700 127.500 16.100 127.600 ;
        RECT 17.500 127.200 17.800 127.900 ;
        RECT 18.300 127.700 20.100 127.900 ;
        RECT 19.400 127.200 19.800 127.400 ;
        RECT 16.200 127.100 17.000 127.200 ;
        RECT 17.400 127.100 18.700 127.200 ;
        RECT 14.000 126.800 14.500 127.100 ;
        RECT 15.900 127.000 18.700 127.100 ;
        RECT 7.800 125.400 8.200 126.200 ;
        RECT 8.600 126.100 9.000 126.200 ;
        RECT 9.400 126.100 9.800 126.200 ;
        RECT 11.000 126.100 11.400 126.200 ;
        RECT 11.800 126.100 12.100 126.800 ;
        RECT 14.200 126.200 14.500 126.800 ;
        RECT 14.800 126.800 18.700 127.000 ;
        RECT 19.400 126.900 20.200 127.200 ;
        RECT 19.800 126.800 20.200 126.900 ;
        RECT 14.800 126.700 16.200 126.800 ;
        RECT 14.800 126.600 15.200 126.700 ;
        RECT 16.600 126.200 16.900 126.800 ;
        RECT 8.600 125.800 9.800 126.100 ;
        RECT 10.600 125.800 12.100 126.100 ;
        RECT 13.400 126.100 13.800 126.200 ;
        RECT 14.200 126.100 14.600 126.200 ;
        RECT 15.500 126.100 15.900 126.200 ;
        RECT 13.400 125.800 14.600 126.100 ;
        RECT 15.100 125.800 15.900 126.100 ;
        RECT 16.600 125.800 17.000 126.200 ;
        RECT 8.700 125.100 9.000 125.800 ;
        RECT 10.600 125.600 11.000 125.800 ;
        RECT 14.200 125.100 14.500 125.800 ;
        RECT 15.100 125.700 15.500 125.800 ;
        RECT 17.400 125.100 17.800 125.200 ;
        RECT 18.400 125.100 18.700 126.800 ;
        RECT 19.000 126.100 19.400 126.600 ;
        RECT 20.600 126.100 21.000 129.900 ;
        RECT 22.200 127.100 22.600 129.900 ;
        RECT 23.800 127.900 24.200 129.900 ;
        RECT 26.000 128.100 26.800 129.900 ;
        RECT 23.800 127.600 25.000 127.900 ;
        RECT 24.600 127.500 25.000 127.600 ;
        RECT 25.300 127.400 25.700 127.800 ;
        RECT 25.300 127.200 25.600 127.400 ;
        RECT 19.000 125.800 21.000 126.100 ;
        RECT 21.400 126.800 22.600 127.100 ;
        RECT 25.200 126.800 25.600 127.200 ;
        RECT 26.000 127.100 26.300 128.100 ;
        RECT 28.600 127.900 29.000 129.900 ;
        RECT 29.700 129.200 30.100 129.900 ;
        RECT 29.400 128.800 30.100 129.200 ;
        RECT 29.700 128.200 30.100 128.800 ;
        RECT 29.700 127.900 30.600 128.200 ;
        RECT 26.600 127.400 27.400 127.800 ;
        RECT 27.700 127.600 29.000 127.900 ;
        RECT 27.700 127.500 28.100 127.600 ;
        RECT 26.000 126.800 26.500 127.100 ;
        RECT 21.400 126.200 21.700 126.800 ;
        RECT 21.400 125.800 21.800 126.200 ;
        RECT 3.800 121.100 4.200 123.100 ;
        RECT 5.400 121.100 5.800 125.100 ;
        RECT 7.000 124.700 7.900 125.100 ;
        RECT 7.500 121.100 7.900 124.700 ;
        RECT 8.600 121.100 9.000 125.100 ;
        RECT 9.400 124.800 11.400 125.100 ;
        RECT 9.400 121.100 9.800 124.800 ;
        RECT 11.000 121.100 11.400 124.800 ;
        RECT 11.800 124.800 13.000 125.100 ;
        RECT 11.800 121.100 12.200 124.800 ;
        RECT 12.600 124.700 13.000 124.800 ;
        RECT 14.000 121.100 14.800 125.100 ;
        RECT 15.700 124.800 17.000 125.100 ;
        RECT 17.400 124.800 18.100 125.100 ;
        RECT 18.400 124.800 18.900 125.100 ;
        RECT 15.700 124.700 16.100 124.800 ;
        RECT 16.600 121.100 17.000 124.800 ;
        RECT 17.800 124.200 18.100 124.800 ;
        RECT 17.800 123.800 18.200 124.200 ;
        RECT 18.500 121.100 18.900 124.800 ;
        RECT 20.600 121.100 21.000 125.800 ;
        RECT 22.200 121.100 22.600 126.800 ;
        RECT 26.200 126.200 26.500 126.800 ;
        RECT 26.200 125.800 26.600 126.200 ;
        RECT 27.500 126.100 27.900 126.200 ;
        RECT 27.100 125.800 27.900 126.100 ;
        RECT 26.200 125.200 26.500 125.800 ;
        RECT 27.100 125.700 27.500 125.800 ;
        RECT 26.200 125.100 27.400 125.200 ;
        RECT 23.800 124.800 25.000 125.100 ;
        RECT 23.800 121.100 24.200 124.800 ;
        RECT 24.600 124.700 25.000 124.800 ;
        RECT 26.000 124.800 27.400 125.100 ;
        RECT 27.700 124.800 29.000 125.100 ;
        RECT 26.000 121.100 26.800 124.800 ;
        RECT 27.700 124.700 28.100 124.800 ;
        RECT 28.600 121.100 29.000 124.800 ;
        RECT 29.400 124.400 29.800 125.200 ;
        RECT 30.200 121.100 30.600 127.900 ;
        RECT 31.000 126.800 31.400 127.600 ;
        RECT 31.800 127.500 32.200 129.900 ;
        RECT 34.000 129.200 34.400 129.900 ;
        RECT 33.400 128.900 34.400 129.200 ;
        RECT 36.200 128.900 36.600 129.900 ;
        RECT 38.300 129.200 38.900 129.900 ;
        RECT 38.200 128.900 38.900 129.200 ;
        RECT 33.400 128.500 33.800 128.900 ;
        RECT 36.200 128.600 36.500 128.900 ;
        RECT 34.200 128.200 34.600 128.600 ;
        RECT 35.100 128.300 36.500 128.600 ;
        RECT 38.200 128.500 38.600 128.900 ;
        RECT 35.100 128.200 35.500 128.300 ;
        RECT 32.200 127.100 33.000 127.200 ;
        RECT 34.300 127.100 34.600 128.200 ;
        RECT 39.100 127.700 39.500 127.800 ;
        RECT 40.600 127.700 41.000 129.900 ;
        RECT 39.100 127.400 41.000 127.700 ;
        RECT 35.000 127.100 35.400 127.200 ;
        RECT 37.100 127.100 37.500 127.200 ;
        RECT 32.200 126.800 37.700 127.100 ;
        RECT 33.700 126.700 34.100 126.800 ;
        RECT 32.900 126.200 33.300 126.300 ;
        RECT 34.200 126.200 34.600 126.300 ;
        RECT 37.400 126.200 37.700 126.800 ;
        RECT 38.200 126.400 38.600 126.500 ;
        RECT 32.900 125.900 35.400 126.200 ;
        RECT 35.000 125.800 35.400 125.900 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 38.200 126.100 40.100 126.400 ;
        RECT 39.700 126.000 40.100 126.100 ;
        RECT 31.800 125.500 34.600 125.600 ;
        RECT 31.800 125.400 34.700 125.500 ;
        RECT 31.800 125.300 36.700 125.400 ;
        RECT 31.800 121.100 32.200 125.300 ;
        RECT 34.300 125.100 36.700 125.300 ;
        RECT 33.400 124.500 36.100 124.800 ;
        RECT 33.400 124.400 33.800 124.500 ;
        RECT 35.700 124.400 36.100 124.500 ;
        RECT 36.400 124.500 36.700 125.100 ;
        RECT 37.400 125.200 37.700 125.800 ;
        RECT 38.900 125.700 39.300 125.800 ;
        RECT 40.600 125.700 41.000 127.400 ;
        RECT 42.200 128.900 42.600 129.900 ;
        RECT 42.200 127.200 42.500 128.900 ;
        RECT 43.000 127.800 43.400 128.600 ;
        RECT 44.100 128.400 44.500 129.900 ;
        RECT 43.800 127.900 44.500 128.400 ;
        RECT 46.200 127.900 46.600 129.900 ;
        RECT 47.800 128.900 48.200 129.900 ;
        RECT 42.200 126.800 42.600 127.200 ;
        RECT 38.900 125.400 41.000 125.700 ;
        RECT 41.400 125.400 41.800 126.200 ;
        RECT 37.400 124.900 38.600 125.200 ;
        RECT 37.100 124.500 37.500 124.600 ;
        RECT 36.400 124.200 37.500 124.500 ;
        RECT 38.300 124.400 38.600 124.900 ;
        RECT 38.300 124.000 39.000 124.400 ;
        RECT 35.100 123.700 35.500 123.800 ;
        RECT 36.500 123.700 36.900 123.800 ;
        RECT 33.400 123.100 33.800 123.500 ;
        RECT 35.100 123.400 36.900 123.700 ;
        RECT 36.200 123.100 36.500 123.400 ;
        RECT 38.200 123.100 38.600 123.500 ;
        RECT 33.400 122.800 34.400 123.100 ;
        RECT 34.000 121.100 34.400 122.800 ;
        RECT 36.200 121.100 36.600 123.100 ;
        RECT 38.300 121.100 38.900 123.100 ;
        RECT 40.600 121.100 41.000 125.400 ;
        RECT 42.200 125.100 42.500 126.800 ;
        RECT 43.800 126.200 44.100 127.900 ;
        RECT 46.200 127.800 46.500 127.900 ;
        RECT 45.600 127.600 46.500 127.800 ;
        RECT 44.400 127.500 46.500 127.600 ;
        RECT 44.400 127.300 45.900 127.500 ;
        RECT 44.400 127.200 44.800 127.300 ;
        RECT 43.800 125.800 44.200 126.200 ;
        RECT 43.800 125.200 44.100 125.800 ;
        RECT 44.500 125.500 44.800 127.200 ;
        RECT 47.800 127.200 48.100 128.900 ;
        RECT 52.300 128.200 52.700 129.900 ;
        RECT 51.800 127.900 52.700 128.200 ;
        RECT 47.800 126.800 48.200 127.200 ;
        RECT 51.000 126.800 51.400 127.600 ;
        RECT 44.500 125.200 45.700 125.500 ;
        RECT 41.700 124.700 42.600 125.100 ;
        RECT 41.700 122.200 42.100 124.700 ;
        RECT 41.700 121.800 42.600 122.200 ;
        RECT 41.700 121.100 42.100 121.800 ;
        RECT 43.800 121.100 44.200 125.200 ;
        RECT 45.400 123.100 45.700 125.200 ;
        RECT 47.800 125.200 48.100 126.800 ;
        RECT 47.800 125.100 48.200 125.200 ;
        RECT 47.300 124.700 48.200 125.100 ;
        RECT 45.400 121.100 45.800 123.100 ;
        RECT 47.300 121.100 47.700 124.700 ;
        RECT 51.800 121.100 52.200 127.900 ;
        RECT 53.400 127.800 53.800 128.600 ;
        RECT 54.200 127.100 54.600 129.900 ;
        RECT 55.000 127.900 55.400 129.900 ;
        RECT 57.200 128.100 58.000 129.900 ;
        RECT 55.000 127.600 56.200 127.900 ;
        RECT 55.800 127.500 56.200 127.600 ;
        RECT 56.500 127.400 56.900 127.800 ;
        RECT 56.500 127.200 56.800 127.400 ;
        RECT 55.000 127.100 55.800 127.200 ;
        RECT 54.200 126.800 55.800 127.100 ;
        RECT 56.400 126.800 56.800 127.200 ;
        RECT 52.600 124.400 53.000 125.200 ;
        RECT 54.200 121.100 54.600 126.800 ;
        RECT 57.200 126.400 57.500 128.100 ;
        RECT 59.800 127.900 60.200 129.900 ;
        RECT 57.800 127.700 58.600 127.800 ;
        RECT 57.800 127.400 58.800 127.700 ;
        RECT 59.100 127.600 60.200 127.900 ;
        RECT 59.100 127.500 59.500 127.600 ;
        RECT 60.600 127.500 61.000 129.900 ;
        RECT 62.800 129.200 63.200 129.900 ;
        RECT 62.200 128.900 63.200 129.200 ;
        RECT 65.000 128.900 65.400 129.900 ;
        RECT 67.100 129.200 67.700 129.900 ;
        RECT 67.000 128.900 67.700 129.200 ;
        RECT 62.200 128.500 62.600 128.900 ;
        RECT 65.000 128.600 65.300 128.900 ;
        RECT 63.000 128.200 63.400 128.600 ;
        RECT 63.900 128.300 65.300 128.600 ;
        RECT 67.000 128.500 67.400 128.900 ;
        RECT 63.900 128.200 64.300 128.300 ;
        RECT 58.500 127.200 58.800 127.400 ;
        RECT 57.800 126.700 58.200 127.100 ;
        RECT 58.500 126.900 60.200 127.200 ;
        RECT 59.400 126.800 60.200 126.900 ;
        RECT 61.000 127.100 61.800 127.200 ;
        RECT 63.100 127.100 63.400 128.200 ;
        RECT 67.900 127.700 68.300 127.800 ;
        RECT 69.400 127.700 69.800 129.900 ;
        RECT 67.900 127.400 69.800 127.700 ;
        RECT 70.200 127.900 70.600 129.900 ;
        RECT 72.400 128.100 73.200 129.900 ;
        RECT 70.200 127.600 71.400 127.900 ;
        RECT 71.000 127.500 71.400 127.600 ;
        RECT 65.900 127.100 66.300 127.200 ;
        RECT 61.000 126.800 66.500 127.100 ;
        RECT 62.500 126.700 62.900 126.800 ;
        RECT 57.000 126.200 57.500 126.400 ;
        RECT 56.600 126.100 57.500 126.200 ;
        RECT 57.900 126.400 58.200 126.700 ;
        RECT 57.900 126.100 59.200 126.400 ;
        RECT 56.600 125.800 57.300 126.100 ;
        RECT 58.800 126.000 59.200 126.100 ;
        RECT 61.700 126.200 62.100 126.300 ;
        RECT 63.000 126.200 63.400 126.300 ;
        RECT 66.200 126.200 66.500 126.800 ;
        RECT 67.000 126.400 67.400 126.500 ;
        RECT 61.700 125.900 64.200 126.200 ;
        RECT 63.800 125.800 64.200 125.900 ;
        RECT 66.200 125.800 66.600 126.200 ;
        RECT 67.000 126.100 68.900 126.400 ;
        RECT 68.500 126.000 68.900 126.100 ;
        RECT 57.000 125.100 57.300 125.800 ;
        RECT 57.700 125.700 58.100 125.800 ;
        RECT 57.700 125.400 59.400 125.700 ;
        RECT 59.100 125.100 59.400 125.400 ;
        RECT 60.600 125.500 63.400 125.600 ;
        RECT 60.600 125.400 63.500 125.500 ;
        RECT 60.600 125.300 65.500 125.400 ;
        RECT 55.000 124.800 56.200 125.100 ;
        RECT 57.000 124.800 58.000 125.100 ;
        RECT 55.000 121.100 55.400 124.800 ;
        RECT 55.800 124.700 56.200 124.800 ;
        RECT 57.200 124.200 58.000 124.800 ;
        RECT 59.100 124.800 60.200 125.100 ;
        RECT 59.100 124.700 59.500 124.800 ;
        RECT 57.200 123.800 58.600 124.200 ;
        RECT 57.200 121.100 58.000 123.800 ;
        RECT 59.800 121.100 60.200 124.800 ;
        RECT 60.600 121.100 61.000 125.300 ;
        RECT 63.100 125.100 65.500 125.300 ;
        RECT 62.200 124.500 64.900 124.800 ;
        RECT 62.200 124.400 62.600 124.500 ;
        RECT 64.500 124.400 64.900 124.500 ;
        RECT 65.200 124.500 65.500 125.100 ;
        RECT 66.200 125.200 66.500 125.800 ;
        RECT 67.700 125.700 68.100 125.800 ;
        RECT 69.400 125.700 69.800 127.400 ;
        RECT 71.700 127.400 72.100 127.800 ;
        RECT 71.700 127.200 72.000 127.400 ;
        RECT 70.200 126.800 71.000 127.200 ;
        RECT 71.600 126.800 72.000 127.200 ;
        RECT 72.400 126.400 72.700 128.100 ;
        RECT 75.000 127.900 75.400 129.900 ;
        RECT 73.000 127.700 73.800 127.800 ;
        RECT 73.000 127.400 74.000 127.700 ;
        RECT 74.300 127.600 75.400 127.900 ;
        RECT 75.800 127.900 76.200 129.900 ;
        RECT 78.000 128.100 78.800 129.900 ;
        RECT 75.800 127.600 76.900 127.900 ;
        RECT 77.400 127.700 78.200 127.800 ;
        RECT 74.300 127.500 74.700 127.600 ;
        RECT 76.500 127.500 76.900 127.600 ;
        RECT 73.700 127.200 74.000 127.400 ;
        RECT 77.200 127.400 78.200 127.700 ;
        RECT 77.200 127.200 77.500 127.400 ;
        RECT 73.700 127.100 75.400 127.200 ;
        RECT 75.800 127.100 77.500 127.200 ;
        RECT 73.000 126.700 73.400 127.100 ;
        RECT 73.700 126.900 77.500 127.100 ;
        RECT 74.600 126.800 76.600 126.900 ;
        RECT 72.200 126.200 72.700 126.400 ;
        RECT 71.800 126.100 72.700 126.200 ;
        RECT 73.100 126.400 73.400 126.700 ;
        RECT 77.800 126.700 78.200 127.100 ;
        RECT 77.800 126.400 78.100 126.700 ;
        RECT 73.100 126.100 74.400 126.400 ;
        RECT 71.800 125.800 72.500 126.100 ;
        RECT 74.000 126.000 74.400 126.100 ;
        RECT 76.800 126.100 78.100 126.400 ;
        RECT 78.500 126.400 78.800 128.100 ;
        RECT 80.600 127.900 81.000 129.900 ;
        RECT 79.100 127.400 79.500 127.800 ;
        RECT 79.800 127.600 81.000 127.900 ;
        RECT 79.800 127.500 80.200 127.600 ;
        RECT 79.200 127.200 79.500 127.400 ;
        RECT 79.200 126.800 79.600 127.200 ;
        RECT 80.200 126.800 81.000 127.200 ;
        RECT 81.400 126.800 81.800 127.600 ;
        RECT 82.200 127.100 82.600 129.900 ;
        RECT 83.000 127.900 83.400 129.900 ;
        RECT 85.200 128.100 86.000 129.900 ;
        RECT 83.000 127.600 84.200 127.900 ;
        RECT 83.800 127.500 84.200 127.600 ;
        RECT 84.500 127.400 84.900 127.800 ;
        RECT 84.500 127.200 84.800 127.400 ;
        RECT 83.000 127.100 83.800 127.200 ;
        RECT 82.200 126.800 83.800 127.100 ;
        RECT 84.400 126.800 84.800 127.200 ;
        RECT 78.500 126.200 79.000 126.400 ;
        RECT 78.500 126.100 79.400 126.200 ;
        RECT 76.800 126.000 77.200 126.100 ;
        RECT 78.700 125.800 79.400 126.100 ;
        RECT 80.600 126.100 80.900 126.800 ;
        RECT 82.200 126.100 82.600 126.800 ;
        RECT 85.200 126.400 85.500 128.100 ;
        RECT 87.800 127.900 88.200 129.900 ;
        RECT 85.800 127.700 86.600 127.800 ;
        RECT 85.800 127.400 86.800 127.700 ;
        RECT 87.100 127.600 88.200 127.900 ;
        RECT 87.100 127.500 87.500 127.600 ;
        RECT 86.500 127.200 86.800 127.400 ;
        RECT 85.800 126.700 86.200 127.100 ;
        RECT 86.500 126.900 88.200 127.200 ;
        RECT 90.400 127.100 90.800 129.900 ;
        RECT 91.800 127.900 92.200 129.900 ;
        RECT 92.600 128.000 93.000 129.900 ;
        RECT 94.200 128.000 94.600 129.900 ;
        RECT 92.600 127.900 94.600 128.000 ;
        RECT 91.900 127.200 92.200 127.900 ;
        RECT 92.700 127.700 94.500 127.900 ;
        RECT 93.800 127.200 94.200 127.400 ;
        RECT 90.400 126.900 91.300 127.100 ;
        RECT 87.400 126.800 88.200 126.900 ;
        RECT 90.500 126.800 91.300 126.900 ;
        RECT 91.800 126.800 93.100 127.200 ;
        RECT 93.800 126.900 94.600 127.200 ;
        RECT 95.600 127.100 96.000 129.900 ;
        RECT 98.200 127.900 98.600 129.900 ;
        RECT 99.000 128.000 99.400 129.900 ;
        RECT 100.600 128.000 101.000 129.900 ;
        RECT 105.400 128.900 105.800 129.900 ;
        RECT 107.000 129.200 107.400 129.900 ;
        RECT 99.000 127.900 101.000 128.000 ;
        RECT 105.200 128.800 105.800 128.900 ;
        RECT 106.900 128.800 107.400 129.200 ;
        RECT 105.200 128.500 107.200 128.800 ;
        RECT 98.300 127.200 98.600 127.900 ;
        RECT 99.100 127.700 100.900 127.900 ;
        RECT 100.200 127.200 100.600 127.400 ;
        RECT 94.200 126.800 94.600 126.900 ;
        RECT 95.100 126.900 96.000 127.100 ;
        RECT 95.100 126.800 95.900 126.900 ;
        RECT 98.200 126.800 99.500 127.200 ;
        RECT 100.200 126.900 101.000 127.200 ;
        RECT 100.600 126.800 101.000 126.900 ;
        RECT 85.000 126.200 85.500 126.400 ;
        RECT 80.600 125.800 82.600 126.100 ;
        RECT 84.600 126.100 85.500 126.200 ;
        RECT 85.900 126.400 86.200 126.700 ;
        RECT 85.900 126.100 87.200 126.400 ;
        RECT 84.600 125.800 85.300 126.100 ;
        RECT 86.800 126.000 87.200 126.100 ;
        RECT 89.400 125.800 90.200 126.200 ;
        RECT 67.700 125.400 69.800 125.700 ;
        RECT 66.200 124.900 67.400 125.200 ;
        RECT 65.900 124.500 66.300 124.600 ;
        RECT 65.200 124.200 66.300 124.500 ;
        RECT 67.100 124.400 67.400 124.900 ;
        RECT 67.100 124.000 67.800 124.400 ;
        RECT 63.900 123.700 64.300 123.800 ;
        RECT 65.300 123.700 65.700 123.800 ;
        RECT 62.200 123.100 62.600 123.500 ;
        RECT 63.900 123.400 65.700 123.700 ;
        RECT 65.000 123.100 65.300 123.400 ;
        RECT 67.000 123.100 67.400 123.500 ;
        RECT 62.200 122.800 63.200 123.100 ;
        RECT 62.800 121.100 63.200 122.800 ;
        RECT 65.000 121.100 65.400 123.100 ;
        RECT 67.100 121.100 67.700 123.100 ;
        RECT 69.400 121.100 69.800 125.400 ;
        RECT 72.200 125.100 72.500 125.800 ;
        RECT 72.900 125.700 73.300 125.800 ;
        RECT 77.900 125.700 78.300 125.800 ;
        RECT 72.900 125.400 74.600 125.700 ;
        RECT 74.300 125.100 74.600 125.400 ;
        RECT 76.600 125.400 78.300 125.700 ;
        RECT 76.600 125.100 76.900 125.400 ;
        RECT 78.700 125.200 79.000 125.800 ;
        RECT 78.700 125.100 79.400 125.200 ;
        RECT 70.200 124.800 71.400 125.100 ;
        RECT 72.200 124.800 73.200 125.100 ;
        RECT 70.200 121.100 70.600 124.800 ;
        RECT 71.000 124.700 71.400 124.800 ;
        RECT 72.400 123.200 73.200 124.800 ;
        RECT 74.300 124.800 75.400 125.100 ;
        RECT 74.300 124.700 74.700 124.800 ;
        RECT 72.400 122.800 73.800 123.200 ;
        RECT 72.400 121.100 73.200 122.800 ;
        RECT 75.000 121.100 75.400 124.800 ;
        RECT 75.800 124.800 76.900 125.100 ;
        RECT 75.800 121.100 76.200 124.800 ;
        RECT 76.500 124.700 76.900 124.800 ;
        RECT 78.000 124.800 79.400 125.100 ;
        RECT 79.800 124.800 81.000 125.100 ;
        RECT 78.000 121.100 78.800 124.800 ;
        RECT 79.800 124.700 80.200 124.800 ;
        RECT 80.600 121.100 81.000 124.800 ;
        RECT 82.200 121.100 82.600 125.800 ;
        RECT 85.000 125.100 85.300 125.800 ;
        RECT 85.700 125.700 86.100 125.800 ;
        RECT 85.700 125.400 87.400 125.700 ;
        RECT 87.100 125.100 87.400 125.400 ;
        RECT 83.000 124.800 84.200 125.100 ;
        RECT 85.000 124.800 86.000 125.100 ;
        RECT 83.000 121.100 83.400 124.800 ;
        RECT 83.800 124.700 84.200 124.800 ;
        RECT 85.200 124.200 86.000 124.800 ;
        RECT 87.100 124.800 88.200 125.100 ;
        RECT 88.600 124.800 89.000 125.600 ;
        RECT 91.000 125.200 91.300 126.800 ;
        RECT 91.800 126.100 92.200 126.200 ;
        RECT 92.800 126.100 93.100 126.800 ;
        RECT 91.800 125.800 93.100 126.100 ;
        RECT 93.400 125.800 93.800 126.600 ;
        RECT 91.000 124.800 91.400 125.200 ;
        RECT 91.800 125.100 92.200 125.200 ;
        RECT 92.800 125.100 93.100 125.800 ;
        RECT 95.100 125.200 95.400 126.800 ;
        RECT 96.200 125.800 97.000 126.200 ;
        RECT 99.200 126.100 99.500 126.800 ;
        RECT 97.400 125.800 99.500 126.100 ;
        RECT 99.800 126.100 100.200 126.600 ;
        RECT 101.400 126.100 101.800 126.200 ;
        RECT 99.800 125.800 101.800 126.100 ;
        RECT 91.800 124.800 92.500 125.100 ;
        RECT 92.800 124.800 93.300 125.100 ;
        RECT 95.000 124.800 95.400 125.200 ;
        RECT 97.400 124.800 97.800 125.800 ;
        RECT 98.200 125.100 98.600 125.200 ;
        RECT 99.200 125.100 99.500 125.800 ;
        RECT 105.200 125.200 105.500 128.500 ;
        RECT 106.200 128.100 106.600 128.200 ;
        RECT 107.300 128.100 108.200 128.200 ;
        RECT 106.200 127.800 108.200 128.100 ;
        RECT 109.400 128.000 109.800 129.900 ;
        RECT 111.000 128.000 111.400 129.900 ;
        RECT 109.400 127.900 111.400 128.000 ;
        RECT 111.800 127.900 112.200 129.900 ;
        RECT 112.600 127.900 113.000 129.900 ;
        RECT 114.800 128.100 115.600 129.900 ;
        RECT 109.500 127.700 111.300 127.900 ;
        RECT 109.800 127.200 110.200 127.400 ;
        RECT 111.800 127.200 112.100 127.900 ;
        RECT 112.600 127.600 113.800 127.900 ;
        RECT 113.400 127.500 113.800 127.600 ;
        RECT 114.100 127.400 114.500 127.800 ;
        RECT 114.100 127.200 114.400 127.400 ;
        RECT 106.600 127.100 107.400 127.200 ;
        RECT 107.800 127.100 108.200 127.200 ;
        RECT 106.600 126.800 108.200 127.100 ;
        RECT 109.400 126.900 110.200 127.200 ;
        RECT 109.400 126.800 109.800 126.900 ;
        RECT 110.900 126.800 112.200 127.200 ;
        RECT 112.600 126.800 113.400 127.200 ;
        RECT 114.000 126.800 114.400 127.200 ;
        RECT 105.800 126.100 106.600 126.200 ;
        RECT 107.000 126.100 107.400 126.200 ;
        RECT 105.800 125.800 107.400 126.100 ;
        RECT 110.200 125.800 110.600 126.600 ;
        RECT 110.900 126.200 111.200 126.800 ;
        RECT 114.800 126.400 115.100 128.100 ;
        RECT 117.400 127.900 117.800 129.900 ;
        RECT 115.400 127.700 116.200 127.800 ;
        RECT 115.400 127.400 116.400 127.700 ;
        RECT 116.700 127.600 117.800 127.900 ;
        RECT 119.800 127.900 120.200 129.900 ;
        RECT 120.500 128.200 120.900 128.600 ;
        RECT 120.600 128.100 121.000 128.200 ;
        RECT 121.400 128.100 121.800 128.600 ;
        RECT 116.700 127.500 117.100 127.600 ;
        RECT 116.100 127.200 116.400 127.400 ;
        RECT 115.400 126.700 115.800 127.100 ;
        RECT 116.100 126.900 117.800 127.200 ;
        RECT 117.000 126.800 117.800 126.900 ;
        RECT 114.600 126.200 115.100 126.400 ;
        RECT 110.900 125.800 111.400 126.200 ;
        RECT 114.200 126.100 115.100 126.200 ;
        RECT 115.500 126.400 115.800 126.700 ;
        RECT 119.000 126.400 119.400 127.200 ;
        RECT 119.800 127.100 120.100 127.900 ;
        RECT 120.600 127.800 121.800 128.100 ;
        RECT 121.400 127.100 121.800 127.200 ;
        RECT 119.800 126.800 121.800 127.100 ;
        RECT 115.500 126.100 116.800 126.400 ;
        RECT 114.200 125.800 114.900 126.100 ;
        RECT 116.400 126.000 116.800 126.100 ;
        RECT 118.200 126.100 118.600 126.200 ;
        RECT 119.800 126.100 120.100 126.800 ;
        RECT 120.600 126.100 121.000 126.200 ;
        RECT 118.200 125.800 119.000 126.100 ;
        RECT 119.800 125.800 121.000 126.100 ;
        RECT 121.400 126.100 121.800 126.200 ;
        RECT 122.200 126.100 122.600 129.900 ;
        RECT 124.800 127.100 125.200 129.900 ;
        RECT 126.200 127.900 126.600 129.900 ;
        RECT 128.400 128.100 129.200 129.900 ;
        RECT 126.200 127.600 127.400 127.900 ;
        RECT 127.000 127.500 127.400 127.600 ;
        RECT 127.700 127.400 128.100 127.800 ;
        RECT 127.700 127.200 128.000 127.400 ;
        RECT 124.800 126.900 125.700 127.100 ;
        RECT 124.900 126.800 125.700 126.900 ;
        RECT 126.200 126.800 127.000 127.200 ;
        RECT 127.600 126.800 128.000 127.200 ;
        RECT 121.400 125.800 122.600 126.100 ;
        RECT 123.800 125.800 124.600 126.200 ;
        RECT 98.200 124.800 98.900 125.100 ;
        RECT 99.200 124.800 99.700 125.100 ;
        RECT 103.800 124.900 105.500 125.200 ;
        RECT 110.900 125.100 111.200 125.800 ;
        RECT 111.800 125.100 112.200 125.200 ;
        RECT 114.600 125.100 114.900 125.800 ;
        RECT 115.300 125.700 115.700 125.800 ;
        RECT 115.300 125.400 117.000 125.700 ;
        RECT 118.600 125.600 119.000 125.800 ;
        RECT 116.700 125.100 117.000 125.400 ;
        RECT 120.600 125.100 120.900 125.800 ;
        RECT 103.800 124.800 104.200 124.900 ;
        RECT 87.100 124.700 87.500 124.800 ;
        RECT 85.200 123.800 86.600 124.200 ;
        RECT 85.200 121.100 86.000 123.800 ;
        RECT 87.800 121.100 88.200 124.800 ;
        RECT 90.200 123.800 90.600 124.600 ;
        RECT 91.000 123.500 91.300 124.800 ;
        RECT 92.200 124.200 92.500 124.800 ;
        RECT 92.200 123.800 92.600 124.200 ;
        RECT 89.500 123.200 91.300 123.500 ;
        RECT 89.500 123.100 89.800 123.200 ;
        RECT 89.400 121.100 89.800 123.100 ;
        RECT 91.000 123.100 91.300 123.200 ;
        RECT 91.000 121.100 91.400 123.100 ;
        RECT 92.900 121.100 93.300 124.800 ;
        RECT 95.100 123.500 95.400 124.800 ;
        RECT 95.800 123.800 96.200 124.600 ;
        RECT 98.600 124.200 98.900 124.800 ;
        RECT 98.600 123.800 99.000 124.200 ;
        RECT 95.100 123.200 96.900 123.500 ;
        RECT 95.100 123.100 95.400 123.200 ;
        RECT 95.000 121.100 95.400 123.100 ;
        RECT 96.600 123.100 96.900 123.200 ;
        RECT 96.600 121.100 97.000 123.100 ;
        RECT 99.300 121.100 99.700 124.800 ;
        RECT 103.900 124.500 104.200 124.800 ;
        RECT 110.700 124.800 111.200 125.100 ;
        RECT 111.500 124.800 112.200 125.100 ;
        RECT 112.600 124.800 113.800 125.100 ;
        RECT 114.600 124.800 115.600 125.100 ;
        RECT 104.700 124.500 106.500 124.600 ;
        RECT 103.000 121.500 103.400 124.500 ;
        RECT 103.800 121.700 104.200 124.500 ;
        RECT 104.600 124.300 106.500 124.500 ;
        RECT 103.100 121.400 103.400 121.500 ;
        RECT 104.600 121.500 105.000 124.300 ;
        RECT 106.200 124.100 106.500 124.300 ;
        RECT 107.100 124.400 108.900 124.700 ;
        RECT 107.100 124.100 107.400 124.400 ;
        RECT 104.600 121.400 104.900 121.500 ;
        RECT 103.100 121.100 104.900 121.400 ;
        RECT 105.400 121.400 105.800 124.000 ;
        RECT 106.200 121.700 106.600 124.100 ;
        RECT 107.000 121.400 107.400 124.100 ;
        RECT 105.400 121.100 107.400 121.400 ;
        RECT 108.600 124.100 108.900 124.400 ;
        RECT 108.600 121.100 109.000 124.100 ;
        RECT 110.700 121.100 111.100 124.800 ;
        RECT 111.500 124.200 111.800 124.800 ;
        RECT 111.400 123.800 111.800 124.200 ;
        RECT 112.600 121.100 113.000 124.800 ;
        RECT 113.400 124.700 113.800 124.800 ;
        RECT 114.800 122.200 115.600 124.800 ;
        RECT 116.700 124.800 117.800 125.100 ;
        RECT 116.700 124.700 117.100 124.800 ;
        RECT 114.200 121.800 115.600 122.200 ;
        RECT 114.800 121.100 115.600 121.800 ;
        RECT 117.400 121.100 117.800 124.800 ;
        RECT 118.200 124.800 120.200 125.100 ;
        RECT 118.200 121.100 118.600 124.800 ;
        RECT 119.800 121.100 120.200 124.800 ;
        RECT 120.600 121.100 121.000 125.100 ;
        RECT 122.200 121.100 122.600 125.800 ;
        RECT 123.000 124.800 123.400 125.600 ;
        RECT 125.400 125.200 125.700 126.800 ;
        RECT 128.400 126.400 128.700 128.100 ;
        RECT 131.000 127.900 131.400 129.900 ;
        RECT 129.000 127.700 129.800 127.800 ;
        RECT 129.000 127.400 130.000 127.700 ;
        RECT 130.300 127.600 131.400 127.900 ;
        RECT 130.300 127.500 130.700 127.600 ;
        RECT 129.700 127.200 130.000 127.400 ;
        RECT 129.000 126.700 129.400 127.100 ;
        RECT 129.700 126.900 131.400 127.200 ;
        RECT 133.600 127.100 134.000 129.900 ;
        RECT 135.100 128.200 135.500 128.600 ;
        RECT 135.000 127.800 135.400 128.200 ;
        RECT 135.800 127.900 136.200 129.900 ;
        RECT 138.200 128.000 138.600 129.900 ;
        RECT 139.800 128.000 140.200 129.900 ;
        RECT 138.200 127.900 140.200 128.000 ;
        RECT 140.600 127.900 141.000 129.900 ;
        RECT 141.400 127.900 141.800 129.900 ;
        RECT 143.600 128.100 144.400 129.900 ;
        RECT 135.900 127.200 136.200 127.900 ;
        RECT 138.300 127.700 140.100 127.900 ;
        RECT 138.600 127.200 139.000 127.400 ;
        RECT 140.600 127.200 140.900 127.900 ;
        RECT 141.400 127.600 142.600 127.900 ;
        RECT 142.200 127.500 142.600 127.600 ;
        RECT 142.900 127.400 143.300 127.800 ;
        RECT 142.900 127.200 143.200 127.400 ;
        RECT 133.600 126.900 134.500 127.100 ;
        RECT 130.600 126.800 131.400 126.900 ;
        RECT 133.700 126.800 134.500 126.900 ;
        RECT 135.800 126.800 136.200 127.200 ;
        RECT 128.200 126.200 128.700 126.400 ;
        RECT 127.800 126.100 128.700 126.200 ;
        RECT 129.100 126.400 129.400 126.700 ;
        RECT 129.100 126.100 130.400 126.400 ;
        RECT 127.800 125.800 128.500 126.100 ;
        RECT 130.000 126.000 130.400 126.100 ;
        RECT 132.600 125.800 133.400 126.200 ;
        RECT 125.400 124.800 125.800 125.200 ;
        RECT 128.200 125.100 128.500 125.800 ;
        RECT 128.900 125.700 129.300 125.800 ;
        RECT 128.900 125.400 130.600 125.700 ;
        RECT 130.300 125.100 130.600 125.400 ;
        RECT 126.200 124.800 127.400 125.100 ;
        RECT 128.200 124.800 129.200 125.100 ;
        RECT 124.600 123.800 125.000 124.600 ;
        RECT 125.400 123.500 125.700 124.800 ;
        RECT 123.900 123.200 125.700 123.500 ;
        RECT 123.900 123.100 124.200 123.200 ;
        RECT 123.800 121.100 124.200 123.100 ;
        RECT 125.400 123.100 125.700 123.200 ;
        RECT 125.400 121.100 125.800 123.100 ;
        RECT 126.200 121.100 126.600 124.800 ;
        RECT 127.000 124.700 127.400 124.800 ;
        RECT 128.400 124.200 129.200 124.800 ;
        RECT 130.300 124.800 131.400 125.100 ;
        RECT 131.800 124.800 132.200 125.600 ;
        RECT 134.200 125.200 134.500 126.800 ;
        RECT 135.000 126.100 135.400 126.200 ;
        RECT 135.900 126.100 136.200 126.800 ;
        RECT 136.600 126.400 137.000 127.200 ;
        RECT 138.200 126.900 139.000 127.200 ;
        RECT 138.200 126.800 138.600 126.900 ;
        RECT 139.700 126.800 141.000 127.200 ;
        RECT 141.400 126.800 142.200 127.200 ;
        RECT 142.800 126.800 143.200 127.200 ;
        RECT 143.600 127.100 143.900 128.100 ;
        RECT 146.200 127.900 146.600 129.900 ;
        RECT 147.800 128.900 148.200 129.900 ;
        RECT 144.200 127.400 145.000 127.800 ;
        RECT 145.300 127.600 146.600 127.900 ;
        RECT 147.000 127.800 147.400 128.600 ;
        RECT 145.300 127.500 145.700 127.600 ;
        RECT 147.900 127.200 148.200 128.900 ;
        RECT 145.800 127.100 146.600 127.200 ;
        RECT 143.600 126.800 144.100 127.100 ;
        RECT 145.500 127.000 146.600 127.100 ;
        RECT 137.400 126.100 137.800 126.200 ;
        RECT 135.000 125.800 136.200 126.100 ;
        RECT 137.000 125.800 137.800 126.100 ;
        RECT 139.000 125.800 139.400 126.600 ;
        RECT 139.700 126.200 140.000 126.800 ;
        RECT 143.800 126.200 144.100 126.800 ;
        RECT 144.400 126.800 146.600 127.000 ;
        RECT 147.800 126.800 148.200 127.200 ;
        RECT 144.400 126.700 145.800 126.800 ;
        RECT 144.400 126.600 144.800 126.700 ;
        RECT 139.700 125.800 140.200 126.200 ;
        RECT 143.800 126.100 144.200 126.200 ;
        RECT 145.100 126.100 145.500 126.200 ;
        RECT 140.600 125.800 144.200 126.100 ;
        RECT 144.700 125.800 145.500 126.100 ;
        RECT 134.200 124.800 134.600 125.200 ;
        RECT 135.100 125.100 135.400 125.800 ;
        RECT 137.000 125.600 137.400 125.800 ;
        RECT 139.700 125.100 140.000 125.800 ;
        RECT 140.600 125.200 140.900 125.800 ;
        RECT 140.600 125.100 141.000 125.200 ;
        RECT 143.800 125.100 144.100 125.800 ;
        RECT 144.700 125.700 145.100 125.800 ;
        RECT 147.900 125.100 148.200 126.800 ;
        RECT 148.600 126.100 149.000 126.200 ;
        RECT 150.200 126.100 150.600 126.200 ;
        RECT 148.600 125.800 150.600 126.100 ;
        RECT 148.600 125.400 149.000 125.800 ;
        RECT 130.300 124.700 130.700 124.800 ;
        RECT 127.800 123.800 129.200 124.200 ;
        RECT 128.400 121.100 129.200 123.800 ;
        RECT 131.000 121.100 131.400 124.800 ;
        RECT 133.400 123.800 133.800 124.600 ;
        RECT 134.200 123.500 134.500 124.800 ;
        RECT 132.700 123.200 134.500 123.500 ;
        RECT 132.700 123.100 133.000 123.200 ;
        RECT 132.600 121.100 133.000 123.100 ;
        RECT 134.200 121.100 134.600 123.200 ;
        RECT 135.000 121.100 135.400 125.100 ;
        RECT 135.800 124.800 137.800 125.100 ;
        RECT 135.800 121.100 136.200 124.800 ;
        RECT 137.400 121.100 137.800 124.800 ;
        RECT 139.500 124.800 140.000 125.100 ;
        RECT 140.300 124.800 141.000 125.100 ;
        RECT 141.400 124.800 142.600 125.100 ;
        RECT 139.500 121.100 139.900 124.800 ;
        RECT 140.300 124.200 140.600 124.800 ;
        RECT 140.200 123.800 140.600 124.200 ;
        RECT 141.400 121.100 141.800 124.800 ;
        RECT 142.200 124.700 142.600 124.800 ;
        RECT 143.600 121.100 144.400 125.100 ;
        RECT 145.300 124.800 146.600 125.100 ;
        RECT 145.300 124.700 145.700 124.800 ;
        RECT 146.200 121.100 146.600 124.800 ;
        RECT 147.800 124.700 148.700 125.100 ;
        RECT 148.300 122.200 148.700 124.700 ;
        RECT 148.300 121.800 149.000 122.200 ;
        RECT 148.300 121.100 148.700 121.800 ;
        RECT 1.400 113.100 1.800 119.900 ;
        RECT 3.000 116.200 3.400 119.900 ;
        RECT 3.800 116.200 4.200 116.300 ;
        RECT 3.000 115.900 4.200 116.200 ;
        RECT 5.200 115.900 6.000 119.900 ;
        RECT 6.900 116.200 7.300 116.300 ;
        RECT 7.800 116.200 8.200 119.900 ;
        RECT 9.900 116.300 10.300 119.900 ;
        RECT 6.900 115.900 8.200 116.200 ;
        RECT 9.400 115.900 10.300 116.300 ;
        RECT 11.000 116.200 11.400 119.900 ;
        RECT 11.800 116.200 12.200 116.300 ;
        RECT 13.200 116.200 14.000 119.900 ;
        RECT 11.000 115.900 12.200 116.200 ;
        RECT 13.000 115.900 14.000 116.200 ;
        RECT 15.100 116.200 15.500 116.300 ;
        RECT 15.800 116.200 16.200 119.900 ;
        RECT 15.100 115.900 16.200 116.200 ;
        RECT 16.600 116.100 17.000 116.200 ;
        RECT 17.400 116.100 17.800 119.900 ;
        RECT 5.400 115.200 5.700 115.900 ;
        RECT 6.300 115.200 6.700 115.300 ;
        RECT 5.400 114.800 5.800 115.200 ;
        RECT 6.300 114.900 7.100 115.200 ;
        RECT 6.700 114.800 7.100 114.900 ;
        RECT 5.400 114.200 5.700 114.800 ;
        RECT 9.500 114.200 9.800 115.900 ;
        RECT 10.200 114.800 10.600 115.600 ;
        RECT 13.000 115.200 13.300 115.900 ;
        RECT 15.100 115.600 15.400 115.900 ;
        RECT 16.600 115.800 17.800 116.100 ;
        RECT 19.500 116.200 19.900 119.900 ;
        RECT 20.200 116.800 20.600 117.200 ;
        RECT 20.300 116.200 20.600 116.800 ;
        RECT 19.500 115.900 20.000 116.200 ;
        RECT 20.300 115.900 21.000 116.200 ;
        RECT 13.700 115.300 15.400 115.600 ;
        RECT 13.700 115.200 14.100 115.300 ;
        RECT 12.600 114.900 13.300 115.200 ;
        RECT 14.800 114.900 15.200 115.000 ;
        RECT 12.600 114.800 13.500 114.900 ;
        RECT 13.000 114.600 13.500 114.800 ;
        RECT 4.400 113.800 4.800 114.200 ;
        RECT 4.500 113.600 4.800 113.800 ;
        RECT 5.200 113.900 5.700 114.200 ;
        RECT 9.400 114.100 9.800 114.200 ;
        RECT 11.000 114.100 11.800 114.200 ;
        RECT 3.800 113.400 4.200 113.500 ;
        RECT 3.000 113.100 4.200 113.400 ;
        RECT 4.500 113.200 4.900 113.600 ;
        RECT 1.400 112.800 2.300 113.100 ;
        RECT 1.900 112.200 2.300 112.800 ;
        RECT 1.900 111.800 2.600 112.200 ;
        RECT 1.900 111.100 2.300 111.800 ;
        RECT 3.000 111.100 3.400 113.100 ;
        RECT 5.200 112.900 5.500 113.900 ;
        RECT 9.400 113.800 11.800 114.100 ;
        RECT 12.400 113.800 12.800 114.200 ;
        RECT 5.800 113.200 6.600 113.600 ;
        RECT 6.900 113.400 7.300 113.500 ;
        RECT 6.900 113.100 8.200 113.400 ;
        RECT 5.200 112.200 6.000 112.900 ;
        RECT 5.200 111.800 6.600 112.200 ;
        RECT 5.200 111.100 6.000 111.800 ;
        RECT 7.800 111.100 8.200 113.100 ;
        RECT 8.600 112.400 9.000 113.200 ;
        RECT 9.500 112.100 9.800 113.800 ;
        RECT 12.500 113.600 12.800 113.800 ;
        RECT 11.800 113.400 12.200 113.500 ;
        RECT 9.400 111.100 9.800 112.100 ;
        RECT 11.000 113.100 12.200 113.400 ;
        RECT 12.500 113.200 12.900 113.600 ;
        RECT 11.000 111.100 11.400 113.100 ;
        RECT 13.200 112.900 13.500 114.600 ;
        RECT 13.900 114.600 15.200 114.900 ;
        RECT 13.900 114.300 14.200 114.600 ;
        RECT 13.800 113.900 14.200 114.300 ;
        RECT 15.400 114.100 16.200 114.200 ;
        RECT 14.500 113.800 16.200 114.100 ;
        RECT 14.500 113.600 14.800 113.800 ;
        RECT 13.800 113.300 14.800 113.600 ;
        RECT 15.100 113.400 15.500 113.500 ;
        RECT 13.800 113.200 14.600 113.300 ;
        RECT 15.100 113.100 16.200 113.400 ;
        RECT 13.200 111.100 14.000 112.900 ;
        RECT 15.800 111.100 16.200 113.100 ;
        RECT 16.600 112.400 17.000 113.200 ;
        RECT 17.400 111.100 17.800 115.800 ;
        RECT 19.000 114.400 19.400 115.200 ;
        RECT 19.700 115.100 20.000 115.900 ;
        RECT 20.600 115.800 21.000 115.900 ;
        RECT 21.400 115.800 21.800 116.600 ;
        RECT 21.400 115.100 21.700 115.800 ;
        RECT 19.700 114.800 21.700 115.100 ;
        RECT 19.700 114.200 20.000 114.800 ;
        RECT 18.200 114.100 18.600 114.200 ;
        RECT 19.700 114.100 21.000 114.200 ;
        RECT 21.400 114.100 21.800 114.200 ;
        RECT 18.200 113.800 19.000 114.100 ;
        RECT 19.700 113.800 21.800 114.100 ;
        RECT 18.600 113.600 19.000 113.800 ;
        RECT 18.300 113.100 20.100 113.300 ;
        RECT 20.600 113.100 20.900 113.800 ;
        RECT 22.200 113.100 22.600 119.900 ;
        RECT 23.800 116.200 24.200 119.900 ;
        RECT 24.600 116.200 25.000 116.300 ;
        RECT 23.800 115.900 25.000 116.200 ;
        RECT 26.000 116.200 26.800 119.900 ;
        RECT 27.700 116.200 28.100 116.300 ;
        RECT 28.600 116.200 29.000 119.900 ;
        RECT 26.000 115.900 27.400 116.200 ;
        RECT 27.700 115.900 29.000 116.200 ;
        RECT 26.200 115.800 27.400 115.900 ;
        RECT 26.200 115.200 26.500 115.800 ;
        RECT 29.400 115.700 29.800 119.900 ;
        RECT 31.600 118.200 32.000 119.900 ;
        RECT 31.000 117.900 32.000 118.200 ;
        RECT 33.800 117.900 34.200 119.900 ;
        RECT 35.900 117.900 36.500 119.900 ;
        RECT 31.000 117.500 31.400 117.900 ;
        RECT 33.800 117.600 34.100 117.900 ;
        RECT 32.700 117.300 34.500 117.600 ;
        RECT 35.800 117.500 36.200 117.900 ;
        RECT 32.700 117.200 33.100 117.300 ;
        RECT 34.100 117.200 34.500 117.300 ;
        RECT 31.000 116.500 31.400 116.600 ;
        RECT 33.300 116.500 33.700 116.600 ;
        RECT 31.000 116.200 33.700 116.500 ;
        RECT 34.000 116.500 35.100 116.800 ;
        RECT 34.000 115.900 34.300 116.500 ;
        RECT 34.700 116.400 35.100 116.500 ;
        RECT 35.900 116.600 36.600 117.000 ;
        RECT 35.900 116.100 36.200 116.600 ;
        RECT 31.900 115.700 34.300 115.900 ;
        RECT 29.400 115.600 34.300 115.700 ;
        RECT 35.000 115.800 36.200 116.100 ;
        RECT 29.400 115.500 32.300 115.600 ;
        RECT 29.400 115.400 32.200 115.500 ;
        RECT 27.100 115.200 27.500 115.300 ;
        RECT 35.000 115.200 35.300 115.800 ;
        RECT 38.200 115.600 38.600 119.900 ;
        RECT 39.300 116.300 39.700 119.900 ;
        RECT 39.300 115.900 40.200 116.300 ;
        RECT 36.500 115.300 38.600 115.600 ;
        RECT 36.500 115.200 36.900 115.300 ;
        RECT 26.200 114.800 26.600 115.200 ;
        RECT 27.100 114.900 27.900 115.200 ;
        RECT 32.600 115.100 33.000 115.200 ;
        RECT 27.500 114.800 27.900 114.900 ;
        RECT 30.500 114.800 33.000 115.100 ;
        RECT 35.000 114.800 35.400 115.200 ;
        RECT 37.300 114.900 37.700 115.000 ;
        RECT 26.200 114.200 26.500 114.800 ;
        RECT 30.500 114.700 30.900 114.800 ;
        RECT 31.800 114.700 32.200 114.800 ;
        RECT 23.000 114.100 23.400 114.200 ;
        RECT 23.800 114.100 24.600 114.200 ;
        RECT 23.000 113.800 24.600 114.100 ;
        RECT 25.200 113.800 25.600 114.200 ;
        RECT 23.000 113.400 23.400 113.800 ;
        RECT 25.300 113.600 25.600 113.800 ;
        RECT 26.000 113.900 26.500 114.200 ;
        RECT 26.800 114.300 27.200 114.400 ;
        RECT 26.800 114.200 28.200 114.300 ;
        RECT 31.300 114.200 31.700 114.300 ;
        RECT 35.000 114.200 35.300 114.800 ;
        RECT 35.800 114.600 37.700 114.900 ;
        RECT 35.800 114.500 36.200 114.600 ;
        RECT 26.800 114.000 29.000 114.200 ;
        RECT 27.900 113.900 29.000 114.000 ;
        RECT 24.600 113.400 25.000 113.500 ;
        RECT 18.200 113.000 20.200 113.100 ;
        RECT 18.200 111.100 18.600 113.000 ;
        RECT 19.800 111.100 20.200 113.000 ;
        RECT 20.600 111.100 21.000 113.100 ;
        RECT 21.700 112.800 22.600 113.100 ;
        RECT 23.800 113.100 25.000 113.400 ;
        RECT 25.300 113.200 25.700 113.600 ;
        RECT 21.700 112.200 22.100 112.800 ;
        RECT 21.400 111.800 22.100 112.200 ;
        RECT 21.700 111.100 22.100 111.800 ;
        RECT 23.800 111.100 24.200 113.100 ;
        RECT 26.000 112.900 26.300 113.900 ;
        RECT 28.200 113.800 29.000 113.900 ;
        RECT 29.800 113.900 35.300 114.200 ;
        RECT 29.800 113.800 30.600 113.900 ;
        RECT 26.600 113.200 27.400 113.600 ;
        RECT 27.700 113.400 28.100 113.500 ;
        RECT 27.700 113.100 29.000 113.400 ;
        RECT 26.000 111.100 26.800 112.900 ;
        RECT 28.600 111.100 29.000 113.100 ;
        RECT 29.400 111.100 29.800 113.500 ;
        RECT 31.900 112.800 32.200 113.900 ;
        RECT 34.700 113.800 35.100 113.900 ;
        RECT 38.200 113.600 38.600 115.300 ;
        RECT 39.000 114.800 39.400 115.600 ;
        RECT 36.700 113.300 38.600 113.600 ;
        RECT 36.700 113.200 37.100 113.300 ;
        RECT 31.000 112.100 31.400 112.500 ;
        RECT 31.800 112.400 32.200 112.800 ;
        RECT 32.700 112.700 33.100 112.800 ;
        RECT 32.700 112.400 34.100 112.700 ;
        RECT 33.800 112.100 34.100 112.400 ;
        RECT 35.800 112.100 36.200 112.500 ;
        RECT 31.000 111.800 32.000 112.100 ;
        RECT 31.600 111.100 32.000 111.800 ;
        RECT 33.800 111.100 34.200 112.100 ;
        RECT 35.800 111.800 36.500 112.100 ;
        RECT 35.900 111.100 36.500 111.800 ;
        RECT 38.200 111.100 38.600 113.300 ;
        RECT 39.800 114.200 40.100 115.900 ;
        RECT 39.800 113.800 40.200 114.200 ;
        RECT 42.200 114.100 42.600 119.900 ;
        RECT 43.000 114.800 43.400 115.200 ;
        RECT 43.800 115.100 44.200 119.900 ;
        RECT 45.900 119.200 46.300 119.900 ;
        RECT 45.400 118.800 46.300 119.200 ;
        RECT 45.900 116.300 46.300 118.800 ;
        RECT 48.300 116.300 48.700 119.900 ;
        RECT 45.400 115.900 46.300 116.300 ;
        RECT 47.800 115.900 48.700 116.300 ;
        RECT 52.300 116.200 52.700 119.900 ;
        RECT 53.000 116.800 53.400 117.200 ;
        RECT 53.100 116.200 53.400 116.800 ;
        RECT 52.300 115.900 52.800 116.200 ;
        RECT 53.100 115.900 53.800 116.200 ;
        RECT 43.800 114.800 44.900 115.100 ;
        RECT 43.000 114.100 43.300 114.800 ;
        RECT 42.200 113.800 43.300 114.100 ;
        RECT 39.000 113.100 39.400 113.200 ;
        RECT 39.800 113.100 40.100 113.800 ;
        RECT 39.000 112.800 40.100 113.100 ;
        RECT 39.800 112.100 40.100 112.800 ;
        RECT 40.600 113.100 41.000 113.200 ;
        RECT 41.400 113.100 41.800 113.200 ;
        RECT 40.600 112.800 41.800 113.100 ;
        RECT 40.600 112.400 41.000 112.800 ;
        RECT 41.400 112.400 41.800 112.800 ;
        RECT 39.800 111.100 40.200 112.100 ;
        RECT 42.200 111.100 42.600 113.800 ;
        RECT 43.000 112.400 43.400 113.200 ;
        RECT 43.800 111.100 44.200 114.800 ;
        RECT 44.600 114.200 44.900 114.800 ;
        RECT 45.500 114.200 45.800 115.900 ;
        RECT 46.200 115.100 46.600 115.600 ;
        RECT 47.900 115.100 48.200 115.900 ;
        RECT 46.200 114.800 48.200 115.100 ;
        RECT 48.600 115.100 49.000 115.600 ;
        RECT 51.800 115.100 52.200 115.200 ;
        RECT 48.600 114.800 52.200 115.100 ;
        RECT 47.900 114.200 48.200 114.800 ;
        RECT 51.800 114.400 52.200 114.800 ;
        RECT 52.500 115.100 52.800 115.900 ;
        RECT 53.400 115.800 53.800 115.900 ;
        RECT 54.200 115.100 54.600 115.200 ;
        RECT 52.500 114.800 54.600 115.100 ;
        RECT 52.500 114.200 52.800 114.800 ;
        RECT 44.600 113.800 45.000 114.200 ;
        RECT 45.400 113.800 45.800 114.200 ;
        RECT 47.800 113.800 48.200 114.200 ;
        RECT 51.000 114.100 51.400 114.200 ;
        RECT 51.000 113.800 51.800 114.100 ;
        RECT 52.500 113.800 53.800 114.200 ;
        RECT 44.600 112.400 45.000 113.200 ;
        RECT 45.500 112.100 45.800 113.800 ;
        RECT 47.000 112.400 47.400 113.200 ;
        RECT 47.900 112.100 48.200 113.800 ;
        RECT 51.400 113.600 51.800 113.800 ;
        RECT 51.100 113.100 52.900 113.300 ;
        RECT 53.400 113.100 53.700 113.800 ;
        RECT 54.200 113.400 54.600 114.200 ;
        RECT 55.000 113.200 55.400 119.900 ;
        RECT 55.800 115.800 56.200 116.600 ;
        RECT 57.900 116.300 58.300 119.900 ;
        RECT 60.300 116.300 60.700 119.900 ;
        RECT 57.400 115.900 58.300 116.300 ;
        RECT 59.800 115.900 60.700 116.300 ;
        RECT 57.500 114.200 57.800 115.900 ;
        RECT 58.200 114.800 58.600 115.600 ;
        RECT 59.000 115.100 59.400 115.200 ;
        RECT 59.900 115.100 60.200 115.900 ;
        RECT 59.000 114.800 60.200 115.100 ;
        RECT 60.600 115.100 61.000 115.600 ;
        RECT 61.400 115.100 61.800 119.900 ;
        RECT 63.000 115.700 63.400 119.900 ;
        RECT 65.200 118.200 65.600 119.900 ;
        RECT 64.600 117.900 65.600 118.200 ;
        RECT 67.400 117.900 67.800 119.900 ;
        RECT 69.500 117.900 70.100 119.900 ;
        RECT 64.600 117.500 65.000 117.900 ;
        RECT 67.400 117.600 67.700 117.900 ;
        RECT 66.300 117.300 68.100 117.600 ;
        RECT 69.400 117.500 69.800 117.900 ;
        RECT 66.300 117.200 66.700 117.300 ;
        RECT 67.700 117.200 68.100 117.300 ;
        RECT 64.600 116.500 65.000 116.600 ;
        RECT 66.900 116.500 67.300 116.600 ;
        RECT 64.600 116.200 67.300 116.500 ;
        RECT 67.600 116.500 68.700 116.800 ;
        RECT 67.600 115.900 67.900 116.500 ;
        RECT 68.300 116.400 68.700 116.500 ;
        RECT 69.500 116.600 70.200 117.000 ;
        RECT 69.500 116.100 69.800 116.600 ;
        RECT 65.500 115.700 67.900 115.900 ;
        RECT 63.000 115.600 67.900 115.700 ;
        RECT 68.600 115.800 69.800 116.100 ;
        RECT 63.000 115.500 65.900 115.600 ;
        RECT 63.000 115.400 65.800 115.500 ;
        RECT 66.200 115.100 66.600 115.200 ;
        RECT 60.600 114.800 61.800 115.100 ;
        RECT 59.900 114.200 60.200 114.800 ;
        RECT 55.800 113.800 56.200 114.200 ;
        RECT 57.400 113.800 57.800 114.200 ;
        RECT 59.800 113.800 60.200 114.200 ;
        RECT 55.800 113.200 56.100 113.800 ;
        RECT 45.400 111.100 45.800 112.100 ;
        RECT 47.800 111.100 48.200 112.100 ;
        RECT 51.000 113.000 53.000 113.100 ;
        RECT 51.000 111.100 51.400 113.000 ;
        RECT 52.600 111.100 53.000 113.000 ;
        RECT 53.400 111.100 53.800 113.100 ;
        RECT 55.000 112.800 56.100 113.200 ;
        RECT 55.500 111.100 55.900 112.800 ;
        RECT 56.600 112.400 57.000 113.200 ;
        RECT 57.500 113.100 57.800 113.800 ;
        RECT 59.000 113.100 59.400 113.200 ;
        RECT 57.400 112.800 59.400 113.100 ;
        RECT 57.500 112.100 57.800 112.800 ;
        RECT 59.000 112.400 59.400 112.800 ;
        RECT 59.900 112.100 60.200 113.800 ;
        RECT 57.400 111.100 57.800 112.100 ;
        RECT 59.800 111.100 60.200 112.100 ;
        RECT 61.400 111.100 61.800 114.800 ;
        RECT 64.100 114.800 66.600 115.100 ;
        RECT 64.100 114.700 64.500 114.800 ;
        RECT 65.400 114.700 65.800 114.800 ;
        RECT 64.900 114.200 65.300 114.300 ;
        RECT 68.600 114.200 68.900 115.800 ;
        RECT 71.800 115.600 72.200 119.900 ;
        RECT 72.600 116.200 73.000 119.900 ;
        RECT 74.800 119.200 75.600 119.900 ;
        RECT 74.800 118.800 76.200 119.200 ;
        RECT 73.300 116.200 73.700 116.300 ;
        RECT 72.600 115.900 73.700 116.200 ;
        RECT 74.800 116.200 75.600 118.800 ;
        RECT 76.600 116.200 77.000 116.300 ;
        RECT 77.400 116.200 77.800 119.900 ;
        RECT 78.300 119.600 80.100 119.900 ;
        RECT 78.300 119.500 78.600 119.600 ;
        RECT 78.200 116.500 78.600 119.500 ;
        RECT 79.800 119.500 80.100 119.600 ;
        RECT 80.600 119.600 82.600 119.900 ;
        RECT 79.000 116.500 79.400 119.300 ;
        RECT 79.800 116.700 80.200 119.500 ;
        RECT 80.600 117.000 81.000 119.600 ;
        RECT 81.400 116.900 81.800 119.300 ;
        RECT 82.200 116.900 82.600 119.600 ;
        RECT 81.400 116.700 81.700 116.900 ;
        RECT 79.800 116.500 81.700 116.700 ;
        RECT 79.100 116.200 79.400 116.500 ;
        RECT 79.900 116.400 81.700 116.500 ;
        RECT 82.300 116.600 82.600 116.900 ;
        RECT 83.800 116.900 84.200 119.900 ;
        RECT 83.800 116.600 84.100 116.900 ;
        RECT 82.300 116.300 84.100 116.600 ;
        RECT 74.800 115.900 75.800 116.200 ;
        RECT 76.600 115.900 77.800 116.200 ;
        RECT 79.000 116.100 79.400 116.200 ;
        RECT 85.900 116.200 86.300 119.900 ;
        RECT 86.600 116.800 87.000 117.200 ;
        RECT 86.700 116.200 87.000 116.800 ;
        RECT 70.100 115.300 72.200 115.600 ;
        RECT 73.400 115.600 73.700 115.900 ;
        RECT 73.400 115.300 75.100 115.600 ;
        RECT 70.100 115.200 70.500 115.300 ;
        RECT 70.900 114.900 71.300 115.000 ;
        RECT 69.400 114.600 71.300 114.900 ;
        RECT 69.400 114.500 69.800 114.600 ;
        RECT 63.400 113.900 68.900 114.200 ;
        RECT 63.400 113.800 64.200 113.900 ;
        RECT 62.200 112.400 62.600 113.200 ;
        RECT 63.000 111.100 63.400 113.500 ;
        RECT 65.500 112.800 65.800 113.900 ;
        RECT 66.200 113.800 66.600 113.900 ;
        RECT 68.300 113.800 68.700 113.900 ;
        RECT 71.800 113.600 72.200 115.300 ;
        RECT 74.700 115.200 75.100 115.300 ;
        RECT 75.500 115.200 75.800 115.900 ;
        RECT 79.000 115.800 80.700 116.100 ;
        RECT 85.900 115.900 86.400 116.200 ;
        RECT 86.700 115.900 87.400 116.200 ;
        RECT 73.600 114.900 74.000 115.000 ;
        RECT 75.500 114.900 76.200 115.200 ;
        RECT 73.600 114.600 74.900 114.900 ;
        RECT 74.600 114.300 74.900 114.600 ;
        RECT 75.300 114.800 76.200 114.900 ;
        RECT 75.300 114.600 75.800 114.800 ;
        RECT 72.600 114.100 73.400 114.200 ;
        RECT 72.600 113.800 74.300 114.100 ;
        RECT 74.600 113.900 75.000 114.300 ;
        RECT 70.300 113.300 72.200 113.600 ;
        RECT 74.000 113.600 74.300 113.800 ;
        RECT 73.300 113.400 73.700 113.500 ;
        RECT 70.300 113.200 70.700 113.300 ;
        RECT 64.600 112.100 65.000 112.500 ;
        RECT 65.400 112.400 65.800 112.800 ;
        RECT 66.300 112.700 66.700 112.800 ;
        RECT 66.300 112.400 67.700 112.700 ;
        RECT 67.400 112.100 67.700 112.400 ;
        RECT 69.400 112.100 69.800 112.500 ;
        RECT 64.600 111.800 65.600 112.100 ;
        RECT 65.200 111.100 65.600 111.800 ;
        RECT 67.400 111.100 67.800 112.100 ;
        RECT 69.400 111.800 70.100 112.100 ;
        RECT 69.500 111.100 70.100 111.800 ;
        RECT 71.800 111.100 72.200 113.300 ;
        RECT 72.600 113.100 73.700 113.400 ;
        RECT 74.000 113.300 75.000 113.600 ;
        RECT 74.200 113.200 75.000 113.300 ;
        RECT 72.600 111.100 73.000 113.100 ;
        RECT 75.300 112.900 75.600 114.600 ;
        RECT 76.000 113.800 76.400 114.200 ;
        RECT 77.000 114.100 77.800 114.200 ;
        RECT 79.000 114.100 79.400 114.200 ;
        RECT 77.000 113.800 79.400 114.100 ;
        RECT 76.000 113.600 76.300 113.800 ;
        RECT 75.900 113.200 76.300 113.600 ;
        RECT 76.600 113.400 77.000 113.500 ;
        RECT 76.600 113.100 77.800 113.400 ;
        RECT 74.800 111.100 75.600 112.900 ;
        RECT 77.400 111.100 77.800 113.100 ;
        RECT 80.400 112.500 80.700 115.800 ;
        RECT 86.100 115.200 86.400 115.900 ;
        RECT 87.000 115.800 87.400 115.900 ;
        RECT 81.000 115.100 81.800 115.200 ;
        RECT 85.400 115.100 85.800 115.200 ;
        RECT 81.000 114.800 85.800 115.100 ;
        RECT 85.400 114.400 85.800 114.800 ;
        RECT 86.100 114.800 86.600 115.200 ;
        RECT 86.100 114.200 86.400 114.800 ;
        RECT 81.400 113.800 82.600 114.200 ;
        RECT 84.600 114.100 85.000 114.200 ;
        RECT 83.000 113.800 85.400 114.100 ;
        RECT 86.100 113.800 87.400 114.200 ;
        RECT 83.000 113.200 83.300 113.800 ;
        RECT 85.000 113.600 85.400 113.800 ;
        RECT 82.500 112.800 83.400 113.200 ;
        RECT 84.700 113.100 86.500 113.300 ;
        RECT 87.000 113.100 87.300 113.800 ;
        RECT 84.600 113.000 86.600 113.100 ;
        RECT 80.400 112.200 82.400 112.500 ;
        RECT 80.400 112.100 81.000 112.200 ;
        RECT 80.600 111.100 81.000 112.100 ;
        RECT 82.100 112.100 82.400 112.200 ;
        RECT 82.100 111.800 82.600 112.100 ;
        RECT 82.200 111.100 82.600 111.800 ;
        RECT 84.600 111.100 85.000 113.000 ;
        RECT 86.200 111.100 86.600 113.000 ;
        RECT 87.000 111.100 87.400 113.100 ;
        RECT 87.800 111.100 88.200 119.900 ;
        RECT 90.200 117.900 90.600 119.900 ;
        RECT 90.300 117.800 90.600 117.900 ;
        RECT 91.800 117.900 92.200 119.900 ;
        RECT 91.800 117.800 92.100 117.900 ;
        RECT 90.300 117.500 92.100 117.800 ;
        RECT 90.200 117.100 90.600 117.200 ;
        RECT 91.000 117.100 91.400 117.200 ;
        RECT 90.200 116.800 91.400 117.100 ;
        RECT 91.000 116.400 91.400 116.800 ;
        RECT 91.800 116.200 92.100 117.500 ;
        RECT 89.400 115.400 89.800 116.200 ;
        RECT 91.800 115.800 92.200 116.200 ;
        RECT 90.200 114.800 91.000 115.200 ;
        RECT 91.800 114.200 92.100 115.800 ;
        RECT 91.300 114.100 92.100 114.200 ;
        RECT 91.200 113.900 92.100 114.100 ;
        RECT 88.600 112.400 89.000 113.200 ;
        RECT 91.200 111.100 91.600 113.900 ;
        RECT 92.600 112.400 93.000 113.200 ;
        RECT 93.400 111.100 93.800 119.900 ;
        RECT 94.200 117.900 94.600 119.900 ;
        RECT 94.300 117.800 94.600 117.900 ;
        RECT 95.800 117.900 96.200 119.900 ;
        RECT 95.800 117.800 96.100 117.900 ;
        RECT 94.300 117.500 96.100 117.800 ;
        RECT 94.300 116.200 94.600 117.500 ;
        RECT 95.000 116.400 95.400 117.200 ;
        RECT 94.200 115.800 94.600 116.200 ;
        RECT 94.300 114.200 94.600 115.800 ;
        RECT 96.600 115.400 97.000 116.200 ;
        RECT 97.400 115.900 97.800 119.900 ;
        RECT 98.200 116.200 98.600 119.900 ;
        RECT 99.800 116.200 100.200 119.900 ;
        RECT 98.200 115.900 100.200 116.200 ;
        RECT 102.200 116.200 102.600 119.900 ;
        RECT 103.800 116.200 104.200 119.900 ;
        RECT 102.200 115.900 104.200 116.200 ;
        RECT 104.600 115.900 105.000 119.900 ;
        RECT 105.400 116.900 105.800 119.900 ;
        RECT 105.500 116.600 105.800 116.900 ;
        RECT 107.000 119.600 109.000 119.900 ;
        RECT 107.000 116.900 107.400 119.600 ;
        RECT 107.800 116.900 108.200 119.300 ;
        RECT 108.600 117.000 109.000 119.600 ;
        RECT 109.500 119.600 111.300 119.900 ;
        RECT 109.500 119.500 109.800 119.600 ;
        RECT 107.000 116.600 107.300 116.900 ;
        RECT 105.500 116.300 107.300 116.600 ;
        RECT 107.900 116.700 108.200 116.900 ;
        RECT 109.400 116.700 109.800 119.500 ;
        RECT 111.000 119.500 111.300 119.600 ;
        RECT 107.900 116.500 109.800 116.700 ;
        RECT 110.200 116.500 110.600 119.300 ;
        RECT 111.000 116.500 111.400 119.500 ;
        RECT 113.100 118.200 113.500 119.900 ;
        RECT 112.600 117.800 113.500 118.200 ;
        RECT 107.900 116.400 109.700 116.500 ;
        RECT 110.200 116.200 110.500 116.500 ;
        RECT 113.100 116.200 113.500 117.800 ;
        RECT 113.800 116.800 114.200 117.200 ;
        RECT 113.900 116.200 114.200 116.800 ;
        RECT 115.000 116.200 115.400 119.900 ;
        RECT 115.700 116.200 116.100 116.300 ;
        RECT 110.200 116.100 110.600 116.200 ;
        RECT 97.500 115.200 97.800 115.900 ;
        RECT 99.400 115.200 99.800 115.400 ;
        RECT 102.600 115.200 103.000 115.400 ;
        RECT 104.600 115.200 104.900 115.900 ;
        RECT 108.900 115.800 110.600 116.100 ;
        RECT 113.100 115.900 113.600 116.200 ;
        RECT 113.900 115.900 114.600 116.200 ;
        RECT 115.000 115.900 116.100 116.200 ;
        RECT 117.200 116.200 118.000 119.900 ;
        RECT 119.000 116.200 119.400 116.300 ;
        RECT 119.800 116.200 120.200 119.900 ;
        RECT 121.400 117.900 121.800 119.900 ;
        RECT 121.500 117.800 121.800 117.900 ;
        RECT 123.000 117.900 123.400 119.900 ;
        RECT 123.800 117.900 124.200 119.900 ;
        RECT 123.000 117.800 123.300 117.900 ;
        RECT 121.500 117.500 123.300 117.800 ;
        RECT 122.200 116.400 122.600 117.200 ;
        RECT 123.000 116.200 123.300 117.500 ;
        RECT 123.900 117.800 124.200 117.900 ;
        RECT 125.400 117.900 125.800 119.900 ;
        RECT 125.400 117.800 125.700 117.900 ;
        RECT 123.900 117.500 125.700 117.800 ;
        RECT 123.900 116.200 124.200 117.500 ;
        RECT 124.600 116.400 125.000 117.200 ;
        RECT 127.000 116.200 127.400 119.900 ;
        RECT 128.600 116.200 129.000 119.900 ;
        RECT 117.200 115.900 118.200 116.200 ;
        RECT 119.000 115.900 120.200 116.200 ;
        RECT 95.400 114.800 96.200 115.200 ;
        RECT 97.400 114.900 98.600 115.200 ;
        RECT 99.400 115.100 100.200 115.200 ;
        RECT 102.200 115.100 103.000 115.200 ;
        RECT 99.400 114.900 103.000 115.100 ;
        RECT 103.800 114.900 105.000 115.200 ;
        RECT 97.400 114.800 97.800 114.900 ;
        RECT 94.300 114.100 95.100 114.200 ;
        RECT 97.400 114.100 97.800 114.200 ;
        RECT 98.300 114.100 98.600 114.900 ;
        RECT 99.800 114.800 102.600 114.900 ;
        RECT 94.300 113.900 95.200 114.100 ;
        RECT 94.800 111.100 95.200 113.900 ;
        RECT 97.400 113.800 98.600 114.100 ;
        RECT 99.000 114.100 99.400 114.600 ;
        RECT 103.000 114.100 103.400 114.600 ;
        RECT 99.000 113.800 103.400 114.100 ;
        RECT 97.400 112.800 97.800 113.200 ;
        RECT 98.300 113.100 98.600 113.800 ;
        RECT 97.500 112.400 97.900 112.800 ;
        RECT 98.200 111.100 98.600 113.100 ;
        RECT 103.800 113.100 104.100 114.900 ;
        RECT 104.600 114.800 105.000 114.900 ;
        RECT 107.000 115.100 107.400 115.200 ;
        RECT 107.800 115.100 108.600 115.200 ;
        RECT 107.000 114.800 108.600 115.100 ;
        RECT 107.000 113.800 108.200 114.200 ;
        RECT 108.900 114.100 109.200 115.800 ;
        RECT 112.600 114.400 113.000 115.200 ;
        RECT 113.300 114.200 113.600 115.900 ;
        RECT 114.200 115.800 114.600 115.900 ;
        RECT 115.800 115.600 116.100 115.900 ;
        RECT 115.800 115.300 117.500 115.600 ;
        RECT 117.100 115.200 117.500 115.300 ;
        RECT 117.900 115.200 118.200 115.900 ;
        RECT 117.900 115.100 118.600 115.200 ;
        RECT 120.600 115.100 121.000 116.200 ;
        RECT 123.000 115.800 123.400 116.200 ;
        RECT 123.800 115.800 124.200 116.200 ;
        RECT 116.000 114.900 116.400 115.000 ;
        RECT 117.900 114.900 121.000 115.100 ;
        RECT 116.000 114.600 117.300 114.900 ;
        RECT 117.000 114.300 117.300 114.600 ;
        RECT 117.700 114.800 121.000 114.900 ;
        RECT 121.400 114.800 122.200 115.200 ;
        RECT 117.700 114.600 118.200 114.800 ;
        RECT 111.800 114.100 112.200 114.200 ;
        RECT 108.900 113.800 112.600 114.100 ;
        RECT 113.300 113.800 114.600 114.200 ;
        RECT 115.000 114.100 115.800 114.200 ;
        RECT 115.000 113.800 116.700 114.100 ;
        RECT 117.000 113.900 117.400 114.300 ;
        RECT 103.800 111.100 104.200 113.100 ;
        RECT 104.600 112.800 105.000 113.200 ;
        RECT 106.200 112.800 107.100 113.200 ;
        RECT 104.500 112.400 104.900 112.800 ;
        RECT 108.900 112.500 109.200 113.800 ;
        RECT 112.200 113.600 112.600 113.800 ;
        RECT 111.900 113.100 113.700 113.300 ;
        RECT 114.200 113.100 114.500 113.800 ;
        RECT 116.400 113.600 116.700 113.800 ;
        RECT 115.700 113.400 116.100 113.500 ;
        RECT 115.000 113.100 116.100 113.400 ;
        RECT 116.400 113.300 117.400 113.600 ;
        RECT 116.600 113.200 117.400 113.300 ;
        RECT 107.200 112.200 109.200 112.500 ;
        RECT 107.200 112.100 107.500 112.200 ;
        RECT 107.000 111.800 107.500 112.100 ;
        RECT 108.600 112.100 109.200 112.200 ;
        RECT 111.800 113.000 113.800 113.100 ;
        RECT 107.000 111.100 107.400 111.800 ;
        RECT 108.600 111.100 109.000 112.100 ;
        RECT 111.800 111.100 112.200 113.000 ;
        RECT 113.400 111.100 113.800 113.000 ;
        RECT 114.200 111.100 114.600 113.100 ;
        RECT 115.000 111.100 115.400 113.100 ;
        RECT 117.700 112.900 118.000 114.600 ;
        RECT 123.000 114.200 123.300 115.800 ;
        RECT 118.400 113.800 118.800 114.200 ;
        RECT 119.400 113.800 120.200 114.200 ;
        RECT 122.500 114.100 123.300 114.200 ;
        RECT 122.400 113.900 123.300 114.100 ;
        RECT 123.900 114.200 124.200 115.800 ;
        RECT 125.000 114.800 125.800 115.200 ;
        RECT 126.200 115.100 126.600 116.200 ;
        RECT 127.000 115.900 129.000 116.200 ;
        RECT 129.400 115.900 129.800 119.900 ;
        RECT 130.200 116.200 130.600 119.900 ;
        RECT 131.000 116.200 131.400 116.300 ;
        RECT 130.200 115.900 131.400 116.200 ;
        RECT 132.400 115.900 133.200 119.900 ;
        RECT 134.100 116.200 134.500 116.300 ;
        RECT 135.000 116.200 135.400 119.900 ;
        RECT 135.800 117.900 136.200 119.900 ;
        RECT 135.900 117.800 136.200 117.900 ;
        RECT 137.400 117.900 137.800 119.900 ;
        RECT 137.400 117.800 137.700 117.900 ;
        RECT 135.900 117.500 137.700 117.800 ;
        RECT 135.900 117.200 136.200 117.500 ;
        RECT 135.800 116.800 136.200 117.200 ;
        RECT 135.900 116.200 136.200 116.800 ;
        RECT 136.600 116.400 137.000 117.200 ;
        RECT 139.000 116.200 139.400 119.900 ;
        RECT 140.600 116.200 141.000 119.900 ;
        RECT 134.100 115.900 135.400 116.200 ;
        RECT 127.400 115.200 127.800 115.400 ;
        RECT 129.400 115.200 129.700 115.900 ;
        RECT 132.600 115.200 132.900 115.900 ;
        RECT 135.800 115.800 136.200 116.200 ;
        RECT 133.500 115.200 133.900 115.300 ;
        RECT 127.000 115.100 127.800 115.200 ;
        RECT 126.200 114.900 127.800 115.100 ;
        RECT 128.600 114.900 129.800 115.200 ;
        RECT 126.200 114.800 127.400 114.900 ;
        RECT 123.900 113.900 125.000 114.200 ;
        RECT 118.400 113.600 118.700 113.800 ;
        RECT 118.300 113.200 118.700 113.600 ;
        RECT 119.000 113.400 119.400 113.500 ;
        RECT 119.000 113.100 120.200 113.400 ;
        RECT 117.200 111.100 118.000 112.900 ;
        RECT 119.800 111.100 120.200 113.100 ;
        RECT 122.400 111.100 122.800 113.900 ;
        RECT 124.400 113.800 125.000 113.900 ;
        RECT 127.800 113.800 128.200 114.600 ;
        RECT 124.400 111.100 124.800 113.800 ;
        RECT 128.600 113.100 128.900 114.900 ;
        RECT 129.400 114.800 129.800 114.900 ;
        RECT 132.600 114.800 133.000 115.200 ;
        RECT 133.500 114.900 134.300 115.200 ;
        RECT 133.900 114.800 134.300 114.900 ;
        RECT 132.600 114.200 132.900 114.800 ;
        RECT 130.200 113.800 131.000 114.200 ;
        RECT 131.600 113.800 132.000 114.200 ;
        RECT 131.700 113.600 132.000 113.800 ;
        RECT 132.400 113.900 132.900 114.200 ;
        RECT 133.200 114.300 133.600 114.400 ;
        RECT 133.200 114.200 134.600 114.300 ;
        RECT 135.900 114.200 136.200 115.800 ;
        RECT 138.200 115.400 138.600 116.200 ;
        RECT 139.000 115.900 141.000 116.200 ;
        RECT 141.400 115.900 141.800 119.900 ;
        RECT 142.200 117.900 142.600 119.900 ;
        RECT 142.300 117.800 142.600 117.900 ;
        RECT 143.800 117.800 144.200 119.900 ;
        RECT 142.300 117.500 144.100 117.800 ;
        RECT 142.300 116.200 142.600 117.500 ;
        RECT 143.000 116.400 143.400 117.200 ;
        RECT 139.400 115.200 139.800 115.400 ;
        RECT 141.400 115.200 141.700 115.900 ;
        RECT 142.200 115.800 142.600 116.200 ;
        RECT 137.000 114.800 137.800 115.200 ;
        RECT 139.000 114.900 139.800 115.200 ;
        RECT 140.600 114.900 141.800 115.200 ;
        RECT 139.000 114.800 139.400 114.900 ;
        RECT 133.200 114.000 135.400 114.200 ;
        RECT 134.300 113.900 135.400 114.000 ;
        RECT 135.900 114.100 136.700 114.200 ;
        RECT 135.900 113.900 136.800 114.100 ;
        RECT 131.000 113.400 131.400 113.500 ;
        RECT 128.600 111.100 129.000 113.100 ;
        RECT 129.400 112.800 129.800 113.200 ;
        RECT 130.200 113.100 131.400 113.400 ;
        RECT 131.700 113.200 132.100 113.600 ;
        RECT 129.300 112.400 129.700 112.800 ;
        RECT 130.200 111.100 130.600 113.100 ;
        RECT 132.400 112.900 132.700 113.900 ;
        RECT 134.600 113.800 135.400 113.900 ;
        RECT 133.000 113.200 133.800 113.600 ;
        RECT 134.100 113.400 134.500 113.500 ;
        RECT 134.100 113.100 135.400 113.400 ;
        RECT 132.400 112.200 133.200 112.900 ;
        RECT 132.400 111.800 133.800 112.200 ;
        RECT 132.400 111.100 133.200 111.800 ;
        RECT 135.000 111.100 135.400 113.100 ;
        RECT 136.400 111.100 136.800 113.900 ;
        RECT 139.800 113.800 140.200 114.600 ;
        RECT 140.600 113.100 140.900 114.900 ;
        RECT 141.400 114.800 141.800 114.900 ;
        RECT 142.300 114.200 142.600 115.800 ;
        RECT 144.600 116.100 145.000 116.200 ;
        RECT 145.400 116.100 145.800 119.900 ;
        RECT 144.600 115.800 145.800 116.100 ;
        RECT 147.000 115.900 147.400 119.900 ;
        RECT 147.800 116.200 148.200 119.900 ;
        RECT 149.400 116.200 149.800 119.900 ;
        RECT 147.800 115.900 149.800 116.200 ;
        RECT 144.600 115.400 145.000 115.800 ;
        RECT 143.400 114.800 144.200 115.200 ;
        RECT 142.300 114.100 143.100 114.200 ;
        RECT 142.300 113.900 143.200 114.100 ;
        RECT 140.600 111.100 141.000 113.100 ;
        RECT 141.400 112.800 141.800 113.200 ;
        RECT 141.300 112.400 141.700 112.800 ;
        RECT 142.800 111.100 143.200 113.900 ;
        RECT 145.400 111.100 145.800 115.800 ;
        RECT 147.100 115.200 147.400 115.900 ;
        RECT 149.000 115.200 149.400 115.400 ;
        RECT 147.000 114.900 148.200 115.200 ;
        RECT 149.000 114.900 149.800 115.200 ;
        RECT 147.000 114.800 147.400 114.900 ;
        RECT 146.200 112.400 146.600 113.200 ;
        RECT 147.000 112.800 147.400 113.200 ;
        RECT 147.900 113.100 148.200 114.900 ;
        RECT 149.400 114.800 149.800 114.900 ;
        RECT 148.600 113.800 149.000 114.600 ;
        RECT 147.100 112.400 147.500 112.800 ;
        RECT 147.800 111.100 148.200 113.100 ;
        RECT 1.400 108.800 1.800 109.900 ;
        RECT 1.500 107.200 1.800 108.800 ;
        RECT 1.400 106.800 1.800 107.200 ;
        RECT 1.500 105.100 1.800 106.800 ;
        RECT 1.400 104.700 2.300 105.100 ;
        RECT 1.900 101.100 2.300 104.700 ;
        RECT 3.800 101.100 4.200 109.900 ;
        RECT 5.400 106.100 5.800 109.900 ;
        RECT 7.000 108.800 7.400 109.900 ;
        RECT 7.000 107.200 7.300 108.800 ;
        RECT 7.800 107.800 8.200 108.600 ;
        RECT 9.900 108.200 10.300 109.900 ;
        RECT 9.400 107.900 10.300 108.200 ;
        RECT 7.000 106.800 7.400 107.200 ;
        RECT 8.600 106.800 9.000 107.600 ;
        RECT 6.200 106.100 6.600 106.200 ;
        RECT 5.400 105.800 6.600 106.100 ;
        RECT 5.400 101.100 5.800 105.800 ;
        RECT 6.200 105.400 6.600 105.800 ;
        RECT 7.000 105.100 7.300 106.800 ;
        RECT 6.500 104.700 7.400 105.100 ;
        RECT 6.500 101.100 6.900 104.700 ;
        RECT 9.400 101.100 9.800 107.900 ;
        RECT 11.000 107.500 11.400 109.900 ;
        RECT 13.200 109.200 13.600 109.900 ;
        RECT 12.600 108.900 13.600 109.200 ;
        RECT 15.400 108.900 15.800 109.900 ;
        RECT 17.500 109.200 18.100 109.900 ;
        RECT 17.400 108.900 18.100 109.200 ;
        RECT 12.600 108.500 13.000 108.900 ;
        RECT 15.400 108.600 15.700 108.900 ;
        RECT 13.400 108.200 13.800 108.600 ;
        RECT 14.300 108.300 15.700 108.600 ;
        RECT 17.400 108.500 17.800 108.900 ;
        RECT 14.300 108.200 14.700 108.300 ;
        RECT 11.400 107.100 12.200 107.200 ;
        RECT 13.500 107.100 13.800 108.200 ;
        RECT 18.300 107.700 18.700 107.800 ;
        RECT 19.800 107.700 20.200 109.900 ;
        RECT 18.300 107.400 20.200 107.700 ;
        RECT 20.600 107.500 21.000 109.900 ;
        RECT 22.800 109.200 23.200 109.900 ;
        RECT 22.200 108.900 23.200 109.200 ;
        RECT 25.000 108.900 25.400 109.900 ;
        RECT 27.100 109.200 27.700 109.900 ;
        RECT 27.000 108.900 27.700 109.200 ;
        RECT 22.200 108.500 22.600 108.900 ;
        RECT 25.000 108.600 25.300 108.900 ;
        RECT 23.000 108.200 23.400 108.600 ;
        RECT 23.900 108.300 25.300 108.600 ;
        RECT 27.000 108.500 27.400 108.900 ;
        RECT 23.900 108.200 24.300 108.300 ;
        RECT 16.300 107.100 16.700 107.200 ;
        RECT 11.400 106.800 16.900 107.100 ;
        RECT 12.900 106.700 13.300 106.800 ;
        RECT 12.100 106.200 12.500 106.300 ;
        RECT 13.400 106.200 13.800 106.300 ;
        RECT 16.600 106.200 16.900 106.800 ;
        RECT 17.400 106.400 17.800 106.500 ;
        RECT 12.100 105.900 14.600 106.200 ;
        RECT 14.200 105.800 14.600 105.900 ;
        RECT 16.600 105.800 17.000 106.200 ;
        RECT 17.400 106.100 19.300 106.400 ;
        RECT 18.900 106.000 19.300 106.100 ;
        RECT 11.000 105.500 13.800 105.600 ;
        RECT 11.000 105.400 13.900 105.500 ;
        RECT 11.000 105.300 15.900 105.400 ;
        RECT 10.200 104.400 10.600 105.200 ;
        RECT 11.000 101.100 11.400 105.300 ;
        RECT 13.500 105.100 15.900 105.300 ;
        RECT 12.600 104.500 15.300 104.800 ;
        RECT 12.600 104.400 13.000 104.500 ;
        RECT 14.900 104.400 15.300 104.500 ;
        RECT 15.600 104.500 15.900 105.100 ;
        RECT 16.600 105.200 16.900 105.800 ;
        RECT 18.100 105.700 18.500 105.800 ;
        RECT 19.800 105.700 20.200 107.400 ;
        RECT 23.100 107.200 23.400 108.200 ;
        RECT 27.900 107.700 28.300 107.800 ;
        RECT 29.400 107.700 29.800 109.900 ;
        RECT 27.900 107.400 29.800 107.700 ;
        RECT 30.200 107.900 30.600 109.900 ;
        RECT 32.400 108.100 33.200 109.900 ;
        RECT 30.200 107.600 31.500 107.900 ;
        RECT 31.100 107.500 31.500 107.600 ;
        RECT 31.800 107.400 32.600 107.800 ;
        RECT 21.000 107.100 21.800 107.200 ;
        RECT 23.000 107.100 23.400 107.200 ;
        RECT 25.900 107.100 26.300 107.200 ;
        RECT 21.000 106.800 26.500 107.100 ;
        RECT 22.500 106.700 22.900 106.800 ;
        RECT 21.700 106.200 22.100 106.300 ;
        RECT 21.700 106.100 24.200 106.200 ;
        RECT 24.600 106.100 25.000 106.200 ;
        RECT 21.700 105.900 25.000 106.100 ;
        RECT 23.800 105.800 25.000 105.900 ;
        RECT 18.100 105.400 20.200 105.700 ;
        RECT 16.600 104.900 17.800 105.200 ;
        RECT 16.300 104.500 16.700 104.600 ;
        RECT 15.600 104.200 16.700 104.500 ;
        RECT 17.500 104.400 17.800 104.900 ;
        RECT 17.500 104.000 18.200 104.400 ;
        RECT 14.300 103.700 14.700 103.800 ;
        RECT 15.700 103.700 16.100 103.800 ;
        RECT 12.600 103.100 13.000 103.500 ;
        RECT 14.300 103.400 16.100 103.700 ;
        RECT 15.400 103.100 15.700 103.400 ;
        RECT 17.400 103.100 17.800 103.500 ;
        RECT 12.600 102.800 13.600 103.100 ;
        RECT 13.200 101.100 13.600 102.800 ;
        RECT 15.400 101.100 15.800 103.100 ;
        RECT 17.500 101.100 18.100 103.100 ;
        RECT 19.800 101.100 20.200 105.400 ;
        RECT 20.600 105.500 23.400 105.600 ;
        RECT 20.600 105.400 23.500 105.500 ;
        RECT 20.600 105.300 25.500 105.400 ;
        RECT 20.600 101.100 21.000 105.300 ;
        RECT 23.100 105.100 25.500 105.300 ;
        RECT 22.200 104.500 24.900 104.800 ;
        RECT 22.200 104.400 22.600 104.500 ;
        RECT 24.500 104.400 24.900 104.500 ;
        RECT 25.200 104.500 25.500 105.100 ;
        RECT 26.200 105.200 26.500 106.800 ;
        RECT 27.000 106.400 27.400 106.500 ;
        RECT 27.000 106.100 28.900 106.400 ;
        RECT 28.500 106.000 28.900 106.100 ;
        RECT 27.700 105.700 28.100 105.800 ;
        RECT 29.400 105.700 29.800 107.400 ;
        RECT 30.200 107.100 31.000 107.200 ;
        RECT 32.900 107.100 33.200 108.100 ;
        RECT 35.000 107.900 35.400 109.900 ;
        RECT 37.100 108.200 37.500 109.900 ;
        RECT 33.500 107.400 33.900 107.800 ;
        RECT 34.200 107.600 35.400 107.900 ;
        RECT 36.600 107.900 37.500 108.200 ;
        RECT 38.200 107.900 38.600 109.900 ;
        RECT 40.400 109.200 41.200 109.900 ;
        RECT 40.400 108.800 41.800 109.200 ;
        RECT 40.400 108.100 41.200 108.800 ;
        RECT 34.200 107.500 34.600 107.600 ;
        RECT 30.200 107.000 31.300 107.100 ;
        RECT 30.200 106.800 32.400 107.000 ;
        RECT 31.000 106.700 32.400 106.800 ;
        RECT 32.000 106.600 32.400 106.700 ;
        RECT 32.700 106.800 33.200 107.100 ;
        RECT 33.600 107.200 33.900 107.400 ;
        RECT 33.600 106.800 34.000 107.200 ;
        RECT 34.600 106.800 35.400 107.200 ;
        RECT 35.800 106.800 36.200 107.600 ;
        RECT 32.700 106.200 33.000 106.800 ;
        RECT 31.300 106.100 31.700 106.200 ;
        RECT 31.300 105.800 32.100 106.100 ;
        RECT 32.600 105.800 33.000 106.200 ;
        RECT 31.700 105.700 32.100 105.800 ;
        RECT 27.700 105.400 29.800 105.700 ;
        RECT 26.200 104.900 27.400 105.200 ;
        RECT 25.900 104.500 26.300 104.600 ;
        RECT 25.200 104.200 26.300 104.500 ;
        RECT 27.100 104.400 27.400 104.900 ;
        RECT 27.100 104.200 27.800 104.400 ;
        RECT 27.100 104.000 28.200 104.200 ;
        RECT 27.500 103.800 28.200 104.000 ;
        RECT 23.900 103.700 24.300 103.800 ;
        RECT 25.300 103.700 25.700 103.800 ;
        RECT 22.200 103.100 22.600 103.500 ;
        RECT 23.900 103.400 25.700 103.700 ;
        RECT 25.000 103.100 25.300 103.400 ;
        RECT 27.000 103.100 27.400 103.500 ;
        RECT 22.200 102.800 23.200 103.100 ;
        RECT 22.800 101.100 23.200 102.800 ;
        RECT 25.000 101.100 25.400 103.100 ;
        RECT 27.100 101.100 27.700 103.100 ;
        RECT 29.400 101.100 29.800 105.400 ;
        RECT 32.700 105.100 33.000 105.800 ;
        RECT 35.800 105.100 36.200 105.200 ;
        RECT 36.600 105.100 37.000 107.900 ;
        RECT 38.200 107.600 39.400 107.900 ;
        RECT 39.000 107.500 39.400 107.600 ;
        RECT 39.700 107.400 40.100 107.800 ;
        RECT 39.700 107.200 40.000 107.400 ;
        RECT 37.400 107.100 37.800 107.200 ;
        RECT 38.200 107.100 39.000 107.200 ;
        RECT 37.400 106.800 39.000 107.100 ;
        RECT 39.600 106.800 40.000 107.200 ;
        RECT 40.400 107.100 40.700 108.100 ;
        RECT 43.000 107.900 43.400 109.900 ;
        RECT 41.000 107.400 41.800 107.800 ;
        RECT 42.100 107.600 43.400 107.900 ;
        RECT 43.800 107.800 44.200 108.600 ;
        RECT 42.100 107.500 42.500 107.600 ;
        RECT 42.600 107.100 43.400 107.200 ;
        RECT 40.400 106.800 40.900 107.100 ;
        RECT 42.300 107.000 43.400 107.100 ;
        RECT 40.600 106.200 40.900 106.800 ;
        RECT 41.200 106.800 43.400 107.000 ;
        RECT 41.200 106.700 42.600 106.800 ;
        RECT 41.200 106.600 41.600 106.700 ;
        RECT 43.000 106.200 43.300 106.800 ;
        RECT 40.600 105.800 41.000 106.200 ;
        RECT 41.900 106.100 42.300 106.200 ;
        RECT 41.500 105.800 42.300 106.100 ;
        RECT 43.000 105.800 43.400 106.200 ;
        RECT 44.600 106.100 45.000 109.900 ;
        RECT 45.400 107.900 45.800 109.900 ;
        RECT 46.200 108.000 46.600 109.900 ;
        RECT 47.800 108.000 48.200 109.900 ;
        RECT 46.200 107.900 48.200 108.000 ;
        RECT 50.200 107.900 50.600 109.900 ;
        RECT 52.400 108.100 53.200 109.900 ;
        RECT 45.500 107.200 45.800 107.900 ;
        RECT 46.300 107.700 48.100 107.900 ;
        RECT 50.200 107.600 51.400 107.900 ;
        RECT 51.000 107.500 51.400 107.600 ;
        RECT 51.700 107.400 52.100 107.800 ;
        RECT 47.400 107.200 47.800 107.400 ;
        RECT 51.700 107.200 52.000 107.400 ;
        RECT 45.400 106.800 46.700 107.200 ;
        RECT 47.400 106.900 48.200 107.200 ;
        RECT 47.800 106.800 48.200 106.900 ;
        RECT 50.200 106.800 51.000 107.200 ;
        RECT 51.600 106.800 52.000 107.200 ;
        RECT 45.400 106.100 45.800 106.200 ;
        RECT 44.600 105.800 45.800 106.100 ;
        RECT 30.200 104.800 31.500 105.100 ;
        RECT 30.200 101.100 30.600 104.800 ;
        RECT 31.100 104.700 31.500 104.800 ;
        RECT 32.400 101.100 33.200 105.100 ;
        RECT 34.200 104.800 35.400 105.100 ;
        RECT 35.800 104.800 37.000 105.100 ;
        RECT 34.200 104.700 34.600 104.800 ;
        RECT 35.000 101.100 35.400 104.800 ;
        RECT 36.600 101.100 37.000 104.800 ;
        RECT 37.400 104.400 37.800 105.200 ;
        RECT 40.600 105.100 40.900 105.800 ;
        RECT 41.500 105.700 41.900 105.800 ;
        RECT 38.200 104.800 39.400 105.100 ;
        RECT 38.200 101.100 38.600 104.800 ;
        RECT 39.000 104.700 39.400 104.800 ;
        RECT 40.400 101.100 41.200 105.100 ;
        RECT 42.100 104.800 43.400 105.100 ;
        RECT 42.100 104.700 42.500 104.800 ;
        RECT 43.000 101.100 43.400 104.800 ;
        RECT 44.600 101.100 45.000 105.800 ;
        RECT 45.400 105.100 45.800 105.200 ;
        RECT 46.400 105.100 46.700 106.800 ;
        RECT 47.000 105.800 47.400 106.600 ;
        RECT 52.400 106.400 52.700 108.100 ;
        RECT 55.000 107.900 55.400 109.900 ;
        RECT 53.000 107.700 53.800 107.800 ;
        RECT 53.000 107.400 54.000 107.700 ;
        RECT 54.300 107.600 55.400 107.900 ;
        RECT 54.300 107.500 54.700 107.600 ;
        RECT 55.800 107.500 56.200 109.900 ;
        RECT 58.000 109.200 58.400 109.900 ;
        RECT 57.400 108.900 58.400 109.200 ;
        RECT 60.200 108.900 60.600 109.900 ;
        RECT 62.300 109.200 62.900 109.900 ;
        RECT 62.200 108.900 62.900 109.200 ;
        RECT 57.400 108.500 57.800 108.900 ;
        RECT 60.200 108.600 60.500 108.900 ;
        RECT 58.200 108.200 58.600 108.600 ;
        RECT 59.100 108.300 60.500 108.600 ;
        RECT 62.200 108.500 62.600 108.900 ;
        RECT 59.100 108.200 59.500 108.300 ;
        RECT 53.700 107.200 54.000 107.400 ;
        RECT 53.000 106.700 53.400 107.100 ;
        RECT 53.700 106.900 55.400 107.200 ;
        RECT 54.600 106.800 55.400 106.900 ;
        RECT 56.200 107.100 57.000 107.200 ;
        RECT 58.300 107.100 58.600 108.200 ;
        RECT 63.100 107.700 63.500 107.800 ;
        RECT 64.600 107.700 65.000 109.900 ;
        RECT 63.100 107.400 65.000 107.700 ;
        RECT 65.400 107.500 65.800 109.900 ;
        RECT 67.600 109.200 68.000 109.900 ;
        RECT 67.000 108.900 68.000 109.200 ;
        RECT 69.800 108.900 70.200 109.900 ;
        RECT 71.900 109.200 72.500 109.900 ;
        RECT 71.800 108.900 72.500 109.200 ;
        RECT 67.000 108.500 67.400 108.900 ;
        RECT 69.800 108.600 70.100 108.900 ;
        RECT 67.800 108.200 68.200 108.600 ;
        RECT 68.700 108.300 70.100 108.600 ;
        RECT 71.800 108.500 72.200 108.900 ;
        RECT 68.700 108.200 69.100 108.300 ;
        RECT 61.100 107.100 61.500 107.200 ;
        RECT 56.200 106.800 61.700 107.100 ;
        RECT 57.700 106.700 58.100 106.800 ;
        RECT 52.200 106.200 52.700 106.400 ;
        RECT 51.800 106.100 52.700 106.200 ;
        RECT 53.100 106.400 53.400 106.700 ;
        RECT 53.100 106.100 54.400 106.400 ;
        RECT 51.800 105.800 52.500 106.100 ;
        RECT 54.000 106.000 54.400 106.100 ;
        RECT 56.900 106.200 57.300 106.300 ;
        RECT 58.200 106.200 58.600 106.300 ;
        RECT 61.400 106.200 61.700 106.800 ;
        RECT 62.200 106.400 62.600 106.500 ;
        RECT 56.900 105.900 59.400 106.200 ;
        RECT 59.000 105.800 59.400 105.900 ;
        RECT 61.400 105.800 61.800 106.200 ;
        RECT 62.200 106.100 64.100 106.400 ;
        RECT 63.700 106.000 64.100 106.100 ;
        RECT 52.200 105.100 52.500 105.800 ;
        RECT 52.900 105.700 53.300 105.800 ;
        RECT 52.900 105.400 54.600 105.700 ;
        RECT 54.300 105.100 54.600 105.400 ;
        RECT 55.800 105.500 58.600 105.600 ;
        RECT 55.800 105.400 58.700 105.500 ;
        RECT 55.800 105.300 60.700 105.400 ;
        RECT 45.400 104.800 46.100 105.100 ;
        RECT 46.400 104.800 46.900 105.100 ;
        RECT 45.800 104.200 46.100 104.800 ;
        RECT 45.800 103.800 46.200 104.200 ;
        RECT 46.500 101.100 46.900 104.800 ;
        RECT 50.200 104.800 51.400 105.100 ;
        RECT 52.200 104.800 53.200 105.100 ;
        RECT 50.200 101.100 50.600 104.800 ;
        RECT 51.000 104.700 51.400 104.800 ;
        RECT 52.400 104.200 53.200 104.800 ;
        RECT 54.300 104.800 55.400 105.100 ;
        RECT 54.300 104.700 54.700 104.800 ;
        RECT 52.400 103.800 53.800 104.200 ;
        RECT 52.400 101.100 53.200 103.800 ;
        RECT 55.000 101.100 55.400 104.800 ;
        RECT 55.800 101.100 56.200 105.300 ;
        RECT 58.300 105.100 60.700 105.300 ;
        RECT 57.400 104.500 60.100 104.800 ;
        RECT 57.400 104.400 57.800 104.500 ;
        RECT 59.700 104.400 60.100 104.500 ;
        RECT 60.400 104.500 60.700 105.100 ;
        RECT 61.400 105.200 61.700 105.800 ;
        RECT 62.900 105.700 63.300 105.800 ;
        RECT 64.600 105.700 65.000 107.400 ;
        RECT 65.800 107.100 66.600 107.200 ;
        RECT 67.900 107.100 68.200 108.200 ;
        RECT 72.700 107.700 73.100 107.800 ;
        RECT 74.200 107.700 74.600 109.900 ;
        RECT 72.700 107.400 74.600 107.700 ;
        RECT 75.000 107.900 75.400 109.900 ;
        RECT 77.200 109.200 78.000 109.900 ;
        RECT 77.200 108.800 78.600 109.200 ;
        RECT 77.200 108.100 78.000 108.800 ;
        RECT 75.000 107.600 76.300 107.900 ;
        RECT 75.900 107.500 76.300 107.600 ;
        RECT 76.600 107.400 77.400 107.800 ;
        RECT 70.700 107.100 71.100 107.200 ;
        RECT 65.800 106.800 71.300 107.100 ;
        RECT 67.300 106.700 67.700 106.800 ;
        RECT 66.500 106.200 66.900 106.300 ;
        RECT 66.500 105.900 69.000 106.200 ;
        RECT 68.600 105.800 69.000 105.900 ;
        RECT 62.900 105.400 65.000 105.700 ;
        RECT 61.400 104.900 62.600 105.200 ;
        RECT 61.100 104.500 61.500 104.600 ;
        RECT 60.400 104.200 61.500 104.500 ;
        RECT 62.300 104.400 62.600 104.900 ;
        RECT 62.300 104.000 63.000 104.400 ;
        RECT 59.100 103.700 59.500 103.800 ;
        RECT 60.500 103.700 60.900 103.800 ;
        RECT 57.400 103.100 57.800 103.500 ;
        RECT 59.100 103.400 60.900 103.700 ;
        RECT 60.200 103.100 60.500 103.400 ;
        RECT 62.200 103.100 62.600 103.500 ;
        RECT 57.400 102.800 58.400 103.100 ;
        RECT 58.000 101.100 58.400 102.800 ;
        RECT 60.200 101.100 60.600 103.100 ;
        RECT 62.300 101.100 62.900 103.100 ;
        RECT 64.600 101.100 65.000 105.400 ;
        RECT 65.400 105.500 68.200 105.600 ;
        RECT 65.400 105.400 68.300 105.500 ;
        RECT 65.400 105.300 70.300 105.400 ;
        RECT 65.400 101.100 65.800 105.300 ;
        RECT 67.900 105.100 70.300 105.300 ;
        RECT 67.000 104.500 69.700 104.800 ;
        RECT 67.000 104.400 67.400 104.500 ;
        RECT 69.300 104.400 69.700 104.500 ;
        RECT 70.000 104.500 70.300 105.100 ;
        RECT 71.000 105.200 71.300 106.800 ;
        RECT 71.800 106.400 72.200 106.500 ;
        RECT 71.800 106.100 73.700 106.400 ;
        RECT 73.300 106.000 73.700 106.100 ;
        RECT 72.500 105.700 72.900 105.800 ;
        RECT 74.200 105.700 74.600 107.400 ;
        RECT 75.000 107.100 75.800 107.200 ;
        RECT 77.700 107.100 78.000 108.100 ;
        RECT 79.800 107.900 80.200 109.900 ;
        RECT 81.900 109.200 82.300 109.900 ;
        RECT 81.400 108.800 82.300 109.200 ;
        RECT 81.900 108.200 82.300 108.800 ;
        RECT 78.300 107.400 78.700 107.800 ;
        RECT 79.000 107.600 80.200 107.900 ;
        RECT 81.400 107.900 82.300 108.200 ;
        RECT 84.600 107.900 85.000 109.900 ;
        RECT 85.300 108.200 85.700 108.600 ;
        RECT 79.000 107.500 79.400 107.600 ;
        RECT 75.000 107.000 76.100 107.100 ;
        RECT 75.000 106.800 77.200 107.000 ;
        RECT 75.800 106.700 77.200 106.800 ;
        RECT 76.800 106.600 77.200 106.700 ;
        RECT 77.500 106.800 78.000 107.100 ;
        RECT 78.400 107.200 78.700 107.400 ;
        RECT 78.400 106.800 78.800 107.200 ;
        RECT 79.400 106.800 80.200 107.200 ;
        RECT 80.600 106.800 81.000 107.600 ;
        RECT 77.500 106.200 77.800 106.800 ;
        RECT 76.100 106.100 76.500 106.200 ;
        RECT 76.100 105.800 76.900 106.100 ;
        RECT 77.400 105.800 77.800 106.200 ;
        RECT 76.500 105.700 76.900 105.800 ;
        RECT 72.500 105.400 74.600 105.700 ;
        RECT 71.000 104.900 72.200 105.200 ;
        RECT 70.700 104.500 71.100 104.600 ;
        RECT 70.000 104.200 71.100 104.500 ;
        RECT 71.900 104.400 72.200 104.900 ;
        RECT 71.900 104.000 72.600 104.400 ;
        RECT 68.700 103.700 69.100 103.800 ;
        RECT 70.100 103.700 70.500 103.800 ;
        RECT 67.000 103.100 67.400 103.500 ;
        RECT 68.700 103.400 70.500 103.700 ;
        RECT 69.800 103.100 70.100 103.400 ;
        RECT 71.800 103.100 72.200 103.500 ;
        RECT 67.000 102.800 68.000 103.100 ;
        RECT 67.600 101.100 68.000 102.800 ;
        RECT 69.800 101.100 70.200 103.100 ;
        RECT 71.900 101.100 72.500 103.100 ;
        RECT 74.200 101.100 74.600 105.400 ;
        RECT 77.500 105.100 77.800 105.800 ;
        RECT 75.000 104.800 76.300 105.100 ;
        RECT 75.000 101.100 75.400 104.800 ;
        RECT 75.900 104.700 76.300 104.800 ;
        RECT 77.200 101.100 78.000 105.100 ;
        RECT 79.000 104.800 80.200 105.100 ;
        RECT 79.000 104.700 79.400 104.800 ;
        RECT 79.800 101.100 80.200 104.800 ;
        RECT 81.400 101.100 81.800 107.900 ;
        RECT 83.800 106.400 84.200 107.200 ;
        RECT 83.000 106.100 83.400 106.200 ;
        RECT 84.600 106.100 84.900 107.900 ;
        RECT 85.400 107.800 85.800 108.200 ;
        RECT 86.800 107.100 87.200 109.900 ;
        RECT 90.000 109.200 90.400 109.900 ;
        RECT 90.000 108.800 90.600 109.200 ;
        RECT 90.000 107.100 90.400 108.800 ;
        RECT 92.700 108.200 93.100 108.600 ;
        RECT 92.600 107.800 93.000 108.200 ;
        RECT 93.400 107.900 93.800 109.900 ;
        RECT 86.300 106.900 87.200 107.100 ;
        RECT 89.500 106.900 90.400 107.100 ;
        RECT 86.300 106.800 87.100 106.900 ;
        RECT 89.500 106.800 90.300 106.900 ;
        RECT 85.400 106.100 85.800 106.200 ;
        RECT 83.000 105.800 83.800 106.100 ;
        RECT 84.600 105.800 85.800 106.100 ;
        RECT 83.400 105.600 83.800 105.800 ;
        RECT 82.200 104.400 82.600 105.200 ;
        RECT 85.400 105.100 85.700 105.800 ;
        RECT 86.300 105.200 86.600 106.800 ;
        RECT 87.400 105.800 88.200 106.200 ;
        RECT 83.000 104.800 85.000 105.100 ;
        RECT 83.000 101.100 83.400 104.800 ;
        RECT 84.600 101.100 85.000 104.800 ;
        RECT 85.400 101.100 85.800 105.100 ;
        RECT 86.200 104.800 86.600 105.200 ;
        RECT 88.600 104.800 89.000 105.600 ;
        RECT 89.500 105.200 89.800 106.800 ;
        RECT 90.600 105.800 91.400 106.200 ;
        RECT 92.600 106.100 93.000 106.200 ;
        RECT 93.500 106.100 93.800 107.900 ;
        RECT 97.400 107.900 97.800 109.900 ;
        RECT 98.100 108.200 98.500 108.600 ;
        RECT 100.300 108.200 100.700 109.900 ;
        RECT 94.200 106.400 94.600 107.200 ;
        RECT 95.000 106.800 95.400 107.200 ;
        RECT 95.000 106.200 95.300 106.800 ;
        RECT 96.600 106.400 97.000 107.200 ;
        RECT 95.000 106.100 95.400 106.200 ;
        RECT 92.600 105.800 93.800 106.100 ;
        RECT 94.600 105.800 95.400 106.100 ;
        RECT 95.800 106.100 96.200 106.200 ;
        RECT 97.400 106.100 97.700 107.900 ;
        RECT 98.200 107.800 98.600 108.200 ;
        RECT 99.800 107.900 100.700 108.200 ;
        RECT 98.200 107.100 98.600 107.200 ;
        RECT 99.000 107.100 99.400 107.600 ;
        RECT 98.200 106.800 99.400 107.100 ;
        RECT 98.200 106.100 98.600 106.200 ;
        RECT 99.000 106.100 99.400 106.200 ;
        RECT 95.800 105.800 96.600 106.100 ;
        RECT 97.400 105.800 99.400 106.100 ;
        RECT 89.400 104.800 89.800 105.200 ;
        RECT 91.800 104.800 92.200 105.600 ;
        RECT 92.700 105.100 93.000 105.800 ;
        RECT 94.600 105.600 95.000 105.800 ;
        RECT 96.200 105.600 96.600 105.800 ;
        RECT 98.200 105.100 98.500 105.800 ;
        RECT 86.300 103.500 86.600 104.800 ;
        RECT 87.000 104.100 87.400 104.600 ;
        RECT 88.600 104.100 89.000 104.200 ;
        RECT 87.000 103.800 89.000 104.100 ;
        RECT 89.500 103.500 89.800 104.800 ;
        RECT 90.200 103.800 90.600 104.600 ;
        RECT 86.300 103.200 88.100 103.500 ;
        RECT 89.500 103.200 91.300 103.500 ;
        RECT 86.300 103.100 86.600 103.200 ;
        RECT 86.200 101.100 86.600 103.100 ;
        RECT 87.800 101.100 88.200 103.200 ;
        RECT 89.500 103.100 89.800 103.200 ;
        RECT 89.400 101.100 89.800 103.100 ;
        RECT 91.000 103.100 91.300 103.200 ;
        RECT 91.000 101.100 91.400 103.100 ;
        RECT 92.600 101.100 93.000 105.100 ;
        RECT 93.400 104.800 95.400 105.100 ;
        RECT 93.400 101.100 93.800 104.800 ;
        RECT 95.000 101.100 95.400 104.800 ;
        RECT 95.800 104.800 97.800 105.100 ;
        RECT 95.800 101.100 96.200 104.800 ;
        RECT 97.400 101.100 97.800 104.800 ;
        RECT 98.200 101.100 98.600 105.100 ;
        RECT 99.800 101.100 100.200 107.900 ;
        RECT 103.600 107.100 104.000 109.900 ;
        RECT 106.800 107.200 107.200 109.900 ;
        RECT 109.400 107.800 109.800 108.600 ;
        RECT 106.800 107.100 107.400 107.200 ;
        RECT 103.100 106.900 104.000 107.100 ;
        RECT 103.100 106.800 103.900 106.900 ;
        RECT 106.300 106.800 107.400 107.100 ;
        RECT 103.100 105.200 103.400 106.800 ;
        RECT 104.200 105.800 105.000 106.200 ;
        RECT 100.600 105.100 101.000 105.200 ;
        RECT 102.200 105.100 102.600 105.200 ;
        RECT 100.600 104.800 102.600 105.100 ;
        RECT 103.000 104.800 103.400 105.200 ;
        RECT 105.400 104.800 105.800 105.600 ;
        RECT 106.300 105.200 106.600 106.800 ;
        RECT 107.400 105.800 108.200 106.200 ;
        RECT 109.400 106.100 109.800 106.200 ;
        RECT 108.600 105.800 109.800 106.100 ;
        RECT 106.200 104.800 106.600 105.200 ;
        RECT 108.600 104.800 109.000 105.800 ;
        RECT 100.600 104.400 101.000 104.800 ;
        RECT 103.100 103.500 103.400 104.800 ;
        RECT 103.800 103.800 104.200 104.600 ;
        RECT 106.300 103.500 106.600 104.800 ;
        RECT 107.000 103.800 107.400 104.600 ;
        RECT 103.100 103.200 104.900 103.500 ;
        RECT 106.300 103.200 108.100 103.500 ;
        RECT 103.100 103.100 103.400 103.200 ;
        RECT 103.000 101.100 103.400 103.100 ;
        RECT 104.600 101.100 105.000 103.200 ;
        RECT 106.300 103.100 106.600 103.200 ;
        RECT 106.200 101.100 106.600 103.100 ;
        RECT 107.800 103.100 108.100 103.200 ;
        RECT 107.800 101.100 108.200 103.100 ;
        RECT 110.200 101.100 110.600 109.900 ;
        RECT 111.000 107.900 111.400 109.900 ;
        RECT 111.800 108.000 112.200 109.900 ;
        RECT 113.400 108.000 113.800 109.900 ;
        RECT 111.800 107.900 113.800 108.000 ;
        RECT 114.200 108.000 114.600 109.900 ;
        RECT 115.800 108.000 116.200 109.900 ;
        RECT 114.200 107.900 116.200 108.000 ;
        RECT 116.600 107.900 117.000 109.900 ;
        RECT 111.100 107.200 111.400 107.900 ;
        RECT 111.900 107.700 113.700 107.900 ;
        RECT 114.300 107.700 116.100 107.900 ;
        RECT 113.000 107.200 113.400 107.400 ;
        RECT 114.600 107.200 115.000 107.400 ;
        RECT 116.600 107.200 116.900 107.900 ;
        RECT 111.000 106.800 112.300 107.200 ;
        RECT 113.000 107.100 113.800 107.200 ;
        RECT 114.200 107.100 115.000 107.200 ;
        RECT 113.000 106.900 115.000 107.100 ;
        RECT 113.400 106.800 114.600 106.900 ;
        RECT 115.700 106.800 117.000 107.200 ;
        RECT 118.000 107.100 118.400 109.900 ;
        RECT 122.200 107.900 122.600 109.900 ;
        RECT 122.900 108.200 123.300 108.600 ;
        RECT 117.500 106.900 118.400 107.100 ;
        RECT 117.500 106.800 118.300 106.900 ;
        RECT 111.000 105.100 111.400 105.200 ;
        RECT 112.000 105.100 112.300 106.800 ;
        RECT 112.600 106.100 113.000 106.600 ;
        RECT 115.000 106.100 115.400 106.600 ;
        RECT 112.600 105.800 115.400 106.100 ;
        RECT 115.700 105.100 116.000 106.800 ;
        RECT 117.500 105.200 117.800 106.800 ;
        RECT 121.400 106.400 121.800 107.200 ;
        RECT 122.200 107.100 122.500 107.900 ;
        RECT 123.000 107.800 123.400 108.200 ;
        RECT 123.800 108.000 124.200 109.900 ;
        RECT 125.400 108.000 125.800 109.900 ;
        RECT 123.800 107.900 125.800 108.000 ;
        RECT 126.200 107.900 126.600 109.900 ;
        RECT 123.900 107.700 125.700 107.900 ;
        RECT 124.200 107.200 124.600 107.400 ;
        RECT 126.200 107.200 126.500 107.900 ;
        RECT 123.800 107.100 124.600 107.200 ;
        RECT 122.200 106.900 124.600 107.100 ;
        RECT 122.200 106.800 124.200 106.900 ;
        RECT 125.300 106.800 126.600 107.200 ;
        RECT 127.600 107.100 128.000 109.900 ;
        RECT 131.800 107.900 132.200 109.900 ;
        RECT 132.500 108.200 132.900 108.600 ;
        RECT 133.500 108.200 133.900 108.600 ;
        RECT 127.100 106.900 128.000 107.100 ;
        RECT 127.100 106.800 127.900 106.900 ;
        RECT 118.600 105.800 119.400 106.200 ;
        RECT 120.600 106.100 121.000 106.200 ;
        RECT 122.200 106.100 122.500 106.800 ;
        RECT 123.000 106.100 123.400 106.200 ;
        RECT 120.600 105.800 121.400 106.100 ;
        RECT 122.200 105.800 123.400 106.100 ;
        RECT 124.600 105.800 125.000 106.600 ;
        RECT 121.000 105.600 121.400 105.800 ;
        RECT 116.600 105.100 117.000 105.200 ;
        RECT 111.000 104.800 111.700 105.100 ;
        RECT 112.000 104.800 112.500 105.100 ;
        RECT 111.400 104.200 111.700 104.800 ;
        RECT 111.400 103.800 111.800 104.200 ;
        RECT 112.100 102.200 112.500 104.800 ;
        RECT 115.500 104.800 116.000 105.100 ;
        RECT 116.300 104.800 117.000 105.100 ;
        RECT 117.400 104.800 117.800 105.200 ;
        RECT 119.800 104.800 120.200 105.600 ;
        RECT 123.000 105.100 123.300 105.800 ;
        RECT 125.300 105.100 125.600 106.800 ;
        RECT 127.100 105.200 127.400 106.800 ;
        RECT 131.000 106.400 131.400 107.200 ;
        RECT 131.800 107.100 132.100 107.900 ;
        RECT 132.600 107.800 133.000 108.200 ;
        RECT 133.400 107.800 133.800 108.200 ;
        RECT 134.200 107.900 134.600 109.900 ;
        RECT 133.400 107.100 133.700 107.800 ;
        RECT 131.800 106.800 133.700 107.100 ;
        RECT 128.200 105.800 129.000 106.200 ;
        RECT 130.200 106.100 130.600 106.200 ;
        RECT 131.800 106.100 132.100 106.800 ;
        RECT 132.600 106.100 133.000 106.200 ;
        RECT 130.200 105.800 131.000 106.100 ;
        RECT 131.800 105.800 133.000 106.100 ;
        RECT 133.400 106.100 133.800 106.200 ;
        RECT 134.300 106.100 134.600 107.900 ;
        RECT 136.600 107.900 137.000 109.900 ;
        RECT 138.800 108.100 139.600 109.900 ;
        RECT 136.600 107.600 137.800 107.900 ;
        RECT 137.400 107.500 137.800 107.600 ;
        RECT 138.100 107.400 138.500 107.800 ;
        RECT 138.100 107.200 138.400 107.400 ;
        RECT 135.000 106.400 135.400 107.200 ;
        RECT 136.600 106.800 137.400 107.200 ;
        RECT 138.000 106.800 138.400 107.200 ;
        RECT 138.800 106.400 139.100 108.100 ;
        RECT 141.400 107.900 141.800 109.900 ;
        RECT 142.200 108.000 142.600 109.900 ;
        RECT 143.800 108.000 144.200 109.900 ;
        RECT 142.200 107.900 144.200 108.000 ;
        RECT 144.600 107.900 145.000 109.900 ;
        RECT 139.400 107.700 140.200 107.800 ;
        RECT 139.400 107.400 140.400 107.700 ;
        RECT 140.700 107.600 141.800 107.900 ;
        RECT 142.300 107.700 144.100 107.900 ;
        RECT 140.700 107.500 141.100 107.600 ;
        RECT 140.100 107.200 140.400 107.400 ;
        RECT 142.600 107.200 143.000 107.400 ;
        RECT 144.600 107.200 144.900 107.900 ;
        RECT 139.400 106.700 139.800 107.100 ;
        RECT 140.100 106.900 141.800 107.200 ;
        RECT 141.000 106.800 141.800 106.900 ;
        RECT 142.200 106.900 143.000 107.200 ;
        RECT 142.200 106.800 142.600 106.900 ;
        RECT 143.700 106.800 145.000 107.200 ;
        RECT 146.000 107.100 146.400 109.900 ;
        RECT 150.200 107.900 150.600 109.900 ;
        RECT 150.900 108.200 151.300 108.600 ;
        RECT 145.500 106.900 146.400 107.100 ;
        RECT 145.500 106.800 146.300 106.900 ;
        RECT 138.600 106.200 139.100 106.400 ;
        RECT 135.800 106.100 136.200 106.200 ;
        RECT 133.400 105.800 134.600 106.100 ;
        RECT 135.400 105.800 136.200 106.100 ;
        RECT 138.200 106.100 139.100 106.200 ;
        RECT 139.500 106.400 139.800 106.700 ;
        RECT 139.500 106.100 140.800 106.400 ;
        RECT 138.200 105.800 138.900 106.100 ;
        RECT 140.400 106.000 140.800 106.100 ;
        RECT 143.000 105.800 143.400 106.600 ;
        RECT 143.700 106.200 144.000 106.800 ;
        RECT 143.700 105.800 144.200 106.200 ;
        RECT 130.600 105.600 131.000 105.800 ;
        RECT 126.200 105.100 126.600 105.200 ;
        RECT 120.600 104.800 122.600 105.100 ;
        RECT 115.500 104.200 115.900 104.800 ;
        RECT 116.300 104.200 116.600 104.800 ;
        RECT 115.000 103.800 115.900 104.200 ;
        RECT 116.200 103.800 116.600 104.200 ;
        RECT 112.100 101.800 113.000 102.200 ;
        RECT 112.100 101.100 112.500 101.800 ;
        RECT 115.500 101.100 115.900 103.800 ;
        RECT 117.500 103.500 117.800 104.800 ;
        RECT 118.200 103.800 118.600 104.600 ;
        RECT 117.500 103.200 119.300 103.500 ;
        RECT 117.500 103.100 117.800 103.200 ;
        RECT 117.400 101.100 117.800 103.100 ;
        RECT 119.000 101.100 119.400 103.200 ;
        RECT 120.600 101.100 121.000 104.800 ;
        RECT 122.200 101.100 122.600 104.800 ;
        RECT 123.000 101.100 123.400 105.100 ;
        RECT 125.100 104.800 125.600 105.100 ;
        RECT 125.900 104.800 126.600 105.100 ;
        RECT 127.000 104.800 127.400 105.200 ;
        RECT 129.400 104.800 129.800 105.600 ;
        RECT 132.600 105.100 132.900 105.800 ;
        RECT 133.500 105.100 133.800 105.800 ;
        RECT 135.400 105.600 135.800 105.800 ;
        RECT 138.600 105.100 138.900 105.800 ;
        RECT 139.300 105.700 139.700 105.800 ;
        RECT 139.300 105.400 141.000 105.700 ;
        RECT 140.700 105.100 141.000 105.400 ;
        RECT 143.700 105.100 144.000 105.800 ;
        RECT 145.500 105.200 145.800 106.800 ;
        RECT 149.400 106.400 149.800 107.200 ;
        RECT 146.600 105.800 147.400 106.200 ;
        RECT 148.600 106.100 149.000 106.200 ;
        RECT 150.200 106.100 150.500 107.900 ;
        RECT 151.000 107.800 151.400 108.200 ;
        RECT 151.000 106.100 151.400 106.200 ;
        RECT 148.600 105.800 149.400 106.100 ;
        RECT 150.200 105.800 151.400 106.100 ;
        RECT 149.000 105.600 149.400 105.800 ;
        RECT 144.600 105.100 145.000 105.200 ;
        RECT 130.200 104.800 132.200 105.100 ;
        RECT 125.100 101.100 125.500 104.800 ;
        RECT 125.900 104.200 126.200 104.800 ;
        RECT 125.800 103.800 126.200 104.200 ;
        RECT 127.100 103.500 127.400 104.800 ;
        RECT 127.800 103.800 128.200 104.600 ;
        RECT 127.100 103.200 128.900 103.500 ;
        RECT 127.100 103.100 127.400 103.200 ;
        RECT 127.000 101.100 127.400 103.100 ;
        RECT 128.600 103.100 128.900 103.200 ;
        RECT 128.600 101.100 129.000 103.100 ;
        RECT 130.200 101.100 130.600 104.800 ;
        RECT 131.800 101.100 132.200 104.800 ;
        RECT 132.600 101.100 133.000 105.100 ;
        RECT 133.400 101.100 133.800 105.100 ;
        RECT 134.200 104.800 136.200 105.100 ;
        RECT 134.200 101.100 134.600 104.800 ;
        RECT 135.800 101.100 136.200 104.800 ;
        RECT 136.600 104.800 137.800 105.100 ;
        RECT 138.600 104.800 139.600 105.100 ;
        RECT 136.600 101.100 137.000 104.800 ;
        RECT 137.400 104.700 137.800 104.800 ;
        RECT 138.800 101.100 139.600 104.800 ;
        RECT 140.700 104.800 141.800 105.100 ;
        RECT 140.700 104.700 141.100 104.800 ;
        RECT 141.400 101.100 141.800 104.800 ;
        RECT 143.500 104.800 144.000 105.100 ;
        RECT 144.300 104.800 145.000 105.100 ;
        RECT 145.400 104.800 145.800 105.200 ;
        RECT 147.800 104.800 148.200 105.600 ;
        RECT 151.000 105.100 151.300 105.800 ;
        RECT 148.600 104.800 150.600 105.100 ;
        RECT 143.500 101.100 143.900 104.800 ;
        RECT 144.300 104.200 144.600 104.800 ;
        RECT 144.200 103.800 144.600 104.200 ;
        RECT 145.500 103.500 145.800 104.800 ;
        RECT 146.200 103.800 146.600 104.600 ;
        RECT 145.500 103.200 147.300 103.500 ;
        RECT 145.500 103.100 145.800 103.200 ;
        RECT 145.400 101.100 145.800 103.100 ;
        RECT 147.000 103.100 147.300 103.200 ;
        RECT 147.000 101.100 147.400 103.100 ;
        RECT 148.600 101.100 149.000 104.800 ;
        RECT 150.200 101.100 150.600 104.800 ;
        RECT 151.000 101.100 151.400 105.100 ;
        RECT 1.400 96.100 1.800 99.900 ;
        RECT 2.200 96.100 2.600 96.600 ;
        RECT 1.400 95.800 2.600 96.100 ;
        RECT 1.400 95.100 1.800 95.800 ;
        RECT 1.400 94.800 2.500 95.100 ;
        RECT 1.400 91.100 1.800 94.800 ;
        RECT 2.200 94.200 2.500 94.800 ;
        RECT 2.200 93.800 2.600 94.200 ;
        RECT 3.000 93.100 3.400 99.900 ;
        RECT 5.900 96.300 6.300 99.900 ;
        RECT 5.400 95.900 6.300 96.300 ;
        RECT 5.500 94.200 5.800 95.900 ;
        RECT 6.200 94.800 6.600 95.600 ;
        RECT 5.400 93.800 5.800 94.200 ;
        RECT 5.500 93.100 5.800 93.800 ;
        RECT 7.800 94.100 8.200 99.900 ;
        RECT 9.400 97.900 9.800 99.900 ;
        RECT 9.500 95.800 9.800 97.900 ;
        RECT 11.000 95.900 11.400 99.900 ;
        RECT 11.800 96.200 12.200 99.900 ;
        RECT 12.600 96.200 13.000 96.300 ;
        RECT 14.000 96.200 14.800 99.900 ;
        RECT 11.800 95.900 13.000 96.200 ;
        RECT 13.800 95.900 14.800 96.200 ;
        RECT 15.900 96.200 16.300 96.300 ;
        RECT 16.600 96.200 17.000 99.900 ;
        RECT 15.900 95.900 17.000 96.200 ;
        RECT 9.500 95.500 10.700 95.800 ;
        RECT 9.400 94.800 9.800 95.200 ;
        RECT 8.600 94.100 9.000 94.600 ;
        RECT 9.500 94.400 9.800 94.800 ;
        RECT 7.800 93.800 9.000 94.100 ;
        RECT 9.400 94.000 10.000 94.400 ;
        RECT 10.400 93.800 10.700 95.500 ;
        RECT 11.100 95.200 11.400 95.900 ;
        RECT 13.800 95.200 14.100 95.900 ;
        RECT 15.900 95.600 16.200 95.900 ;
        RECT 14.500 95.300 16.200 95.600 ;
        RECT 17.400 95.700 17.800 99.900 ;
        RECT 19.600 98.200 20.000 99.900 ;
        RECT 19.000 97.900 20.000 98.200 ;
        RECT 21.800 97.900 22.200 99.900 ;
        RECT 23.900 97.900 24.500 99.900 ;
        RECT 19.000 97.500 19.400 97.900 ;
        RECT 21.800 97.600 22.100 97.900 ;
        RECT 20.700 97.300 22.500 97.600 ;
        RECT 23.800 97.500 24.200 97.900 ;
        RECT 20.700 97.200 21.100 97.300 ;
        RECT 22.100 97.200 22.500 97.300 ;
        RECT 19.000 96.500 19.400 96.600 ;
        RECT 21.300 96.500 21.700 96.600 ;
        RECT 19.000 96.200 21.700 96.500 ;
        RECT 22.000 96.500 23.100 96.800 ;
        RECT 22.000 95.900 22.300 96.500 ;
        RECT 22.700 96.400 23.100 96.500 ;
        RECT 23.900 96.600 24.600 97.000 ;
        RECT 23.900 96.100 24.200 96.600 ;
        RECT 19.900 95.700 22.300 95.900 ;
        RECT 17.400 95.600 22.300 95.700 ;
        RECT 23.000 95.800 24.200 96.100 ;
        RECT 17.400 95.500 20.300 95.600 ;
        RECT 17.400 95.400 20.200 95.500 ;
        RECT 14.500 95.200 14.900 95.300 ;
        RECT 23.000 95.200 23.300 95.800 ;
        RECT 26.200 95.600 26.600 99.900 ;
        RECT 24.500 95.300 26.600 95.600 ;
        RECT 27.000 95.700 27.400 99.900 ;
        RECT 29.200 98.200 29.600 99.900 ;
        RECT 28.600 97.900 29.600 98.200 ;
        RECT 31.400 97.900 31.800 99.900 ;
        RECT 33.500 97.900 34.100 99.900 ;
        RECT 28.600 97.500 29.000 97.900 ;
        RECT 31.400 97.600 31.700 97.900 ;
        RECT 30.300 97.300 32.100 97.600 ;
        RECT 33.400 97.500 33.800 97.900 ;
        RECT 30.300 97.200 30.700 97.300 ;
        RECT 31.700 97.200 32.100 97.300 ;
        RECT 28.600 96.500 29.000 96.600 ;
        RECT 30.900 96.500 31.300 96.600 ;
        RECT 28.600 96.200 31.300 96.500 ;
        RECT 31.600 96.500 32.700 96.800 ;
        RECT 31.600 95.900 31.900 96.500 ;
        RECT 32.300 96.400 32.700 96.500 ;
        RECT 33.500 96.600 34.200 97.000 ;
        RECT 33.500 96.100 33.800 96.600 ;
        RECT 29.500 95.700 31.900 95.900 ;
        RECT 27.000 95.600 31.900 95.700 ;
        RECT 32.600 95.800 33.800 96.100 ;
        RECT 27.000 95.500 29.900 95.600 ;
        RECT 27.000 95.400 29.800 95.500 ;
        RECT 24.500 95.200 24.900 95.300 ;
        RECT 11.000 94.800 11.400 95.200 ;
        RECT 13.400 94.900 14.100 95.200 ;
        RECT 20.600 95.100 21.000 95.200 ;
        RECT 15.600 94.900 16.000 95.000 ;
        RECT 13.400 94.800 14.300 94.900 ;
        RECT 7.000 93.100 7.400 93.200 ;
        RECT 2.500 92.800 3.400 93.100 ;
        RECT 5.400 92.800 7.400 93.100 ;
        RECT 2.500 91.100 2.900 92.800 ;
        RECT 5.500 92.100 5.800 92.800 ;
        RECT 7.000 92.400 7.400 92.800 ;
        RECT 5.400 91.100 5.800 92.100 ;
        RECT 7.800 91.100 8.200 93.800 ;
        RECT 10.400 93.700 10.800 93.800 ;
        RECT 9.300 93.500 10.800 93.700 ;
        RECT 8.700 93.400 10.800 93.500 ;
        RECT 8.700 93.200 9.600 93.400 ;
        RECT 8.700 93.100 9.000 93.200 ;
        RECT 11.100 93.100 11.400 94.800 ;
        RECT 13.800 94.600 14.300 94.800 ;
        RECT 11.800 93.800 12.600 94.200 ;
        RECT 13.200 93.800 13.600 94.200 ;
        RECT 13.300 93.600 13.600 93.800 ;
        RECT 12.600 93.400 13.000 93.500 ;
        RECT 8.600 91.100 9.000 93.100 ;
        RECT 10.700 92.600 11.400 93.100 ;
        RECT 11.800 93.100 13.000 93.400 ;
        RECT 13.300 93.200 13.700 93.600 ;
        RECT 10.700 92.200 11.100 92.600 ;
        RECT 10.700 91.800 11.400 92.200 ;
        RECT 10.700 91.100 11.100 91.800 ;
        RECT 11.800 91.100 12.200 93.100 ;
        RECT 14.000 92.900 14.300 94.600 ;
        RECT 14.700 94.600 16.000 94.900 ;
        RECT 18.500 94.800 21.000 95.100 ;
        RECT 23.000 94.800 23.400 95.200 ;
        RECT 25.300 94.900 25.700 95.000 ;
        RECT 18.500 94.700 18.900 94.800 ;
        RECT 19.800 94.700 20.200 94.800 ;
        RECT 14.700 94.300 15.000 94.600 ;
        RECT 14.600 93.900 15.000 94.300 ;
        RECT 19.300 94.200 19.700 94.300 ;
        RECT 23.000 94.200 23.300 94.800 ;
        RECT 23.800 94.600 25.700 94.900 ;
        RECT 23.800 94.500 24.200 94.600 ;
        RECT 16.200 94.100 17.000 94.200 ;
        RECT 15.300 93.800 17.000 94.100 ;
        RECT 17.800 93.900 23.300 94.200 ;
        RECT 17.800 93.800 18.600 93.900 ;
        RECT 15.300 93.600 15.600 93.800 ;
        RECT 14.600 93.300 15.600 93.600 ;
        RECT 15.900 93.400 16.300 93.500 ;
        RECT 14.600 93.200 15.400 93.300 ;
        RECT 15.900 93.100 17.000 93.400 ;
        RECT 14.000 91.100 14.800 92.900 ;
        RECT 16.600 91.100 17.000 93.100 ;
        RECT 17.400 91.100 17.800 93.500 ;
        RECT 19.900 92.800 20.200 93.900 ;
        RECT 20.600 93.800 21.000 93.900 ;
        RECT 22.700 93.800 23.100 93.900 ;
        RECT 26.200 93.600 26.600 95.300 ;
        RECT 30.200 95.100 30.600 95.200 ;
        RECT 28.100 94.800 30.600 95.100 ;
        RECT 28.100 94.700 28.500 94.800 ;
        RECT 28.900 94.200 29.300 94.300 ;
        RECT 32.600 94.200 32.900 95.800 ;
        RECT 35.800 95.600 36.200 99.900 ;
        RECT 37.900 96.300 38.300 99.900 ;
        RECT 37.400 95.900 38.300 96.300 ;
        RECT 34.100 95.300 36.200 95.600 ;
        RECT 34.100 95.200 34.500 95.300 ;
        RECT 34.900 94.900 35.300 95.000 ;
        RECT 33.400 94.600 35.300 94.900 ;
        RECT 33.400 94.500 33.800 94.600 ;
        RECT 27.400 93.900 32.900 94.200 ;
        RECT 27.400 93.800 28.200 93.900 ;
        RECT 24.700 93.300 26.600 93.600 ;
        RECT 24.700 93.200 25.100 93.300 ;
        RECT 19.000 92.100 19.400 92.500 ;
        RECT 19.800 92.400 20.200 92.800 ;
        RECT 20.700 92.700 21.100 92.800 ;
        RECT 20.700 92.400 22.100 92.700 ;
        RECT 21.800 92.100 22.100 92.400 ;
        RECT 23.800 92.100 24.200 92.500 ;
        RECT 19.000 91.800 20.000 92.100 ;
        RECT 19.600 91.100 20.000 91.800 ;
        RECT 21.800 91.100 22.200 92.100 ;
        RECT 23.800 91.800 24.500 92.100 ;
        RECT 23.900 91.100 24.500 91.800 ;
        RECT 26.200 91.100 26.600 93.300 ;
        RECT 27.000 91.100 27.400 93.500 ;
        RECT 29.500 92.800 29.800 93.900 ;
        RECT 31.000 93.800 31.400 93.900 ;
        RECT 32.300 93.800 32.700 93.900 ;
        RECT 35.800 93.600 36.200 95.300 ;
        RECT 37.500 94.200 37.800 95.900 ;
        RECT 38.200 94.800 38.600 95.600 ;
        RECT 37.400 93.800 37.800 94.200 ;
        RECT 38.200 94.100 38.600 94.200 ;
        RECT 39.000 94.100 39.400 94.200 ;
        RECT 38.200 93.800 39.400 94.100 ;
        RECT 34.300 93.300 36.200 93.600 ;
        RECT 34.300 93.200 34.700 93.300 ;
        RECT 28.600 92.100 29.000 92.500 ;
        RECT 29.400 92.400 29.800 92.800 ;
        RECT 30.300 92.700 30.700 92.800 ;
        RECT 30.300 92.400 31.700 92.700 ;
        RECT 31.400 92.100 31.700 92.400 ;
        RECT 33.400 92.100 33.800 92.500 ;
        RECT 28.600 91.800 29.600 92.100 ;
        RECT 29.200 91.100 29.600 91.800 ;
        RECT 31.400 91.100 31.800 92.100 ;
        RECT 33.400 91.800 34.100 92.100 ;
        RECT 33.500 91.100 34.100 91.800 ;
        RECT 35.800 91.100 36.200 93.300 ;
        RECT 36.600 92.400 37.000 93.200 ;
        RECT 37.500 92.200 37.800 93.800 ;
        RECT 39.000 93.400 39.400 93.800 ;
        RECT 39.800 93.200 40.200 99.900 ;
        RECT 40.600 95.800 41.000 96.600 ;
        RECT 41.400 95.700 41.800 99.900 ;
        RECT 43.600 98.200 44.000 99.900 ;
        RECT 43.000 97.900 44.000 98.200 ;
        RECT 45.800 97.900 46.200 99.900 ;
        RECT 47.900 97.900 48.500 99.900 ;
        RECT 43.000 97.500 43.400 97.900 ;
        RECT 45.800 97.600 46.100 97.900 ;
        RECT 44.700 97.300 46.500 97.600 ;
        RECT 47.800 97.500 48.200 97.900 ;
        RECT 44.700 97.200 45.100 97.300 ;
        RECT 46.100 97.200 46.500 97.300 ;
        RECT 43.000 96.500 43.400 96.600 ;
        RECT 45.300 96.500 45.700 96.600 ;
        RECT 43.000 96.200 45.700 96.500 ;
        RECT 46.000 96.500 47.100 96.800 ;
        RECT 46.000 95.900 46.300 96.500 ;
        RECT 46.700 96.400 47.100 96.500 ;
        RECT 47.900 96.600 48.600 97.000 ;
        RECT 47.900 96.100 48.200 96.600 ;
        RECT 43.900 95.700 46.300 95.900 ;
        RECT 41.400 95.600 46.300 95.700 ;
        RECT 47.000 95.800 48.200 96.100 ;
        RECT 41.400 95.500 44.300 95.600 ;
        RECT 41.400 95.400 44.200 95.500 ;
        RECT 47.000 95.200 47.300 95.800 ;
        RECT 50.200 95.600 50.600 99.900 ;
        RECT 53.900 99.200 54.300 99.900 ;
        RECT 53.900 98.800 54.600 99.200 ;
        RECT 53.900 96.300 54.300 98.800 ;
        RECT 53.400 95.900 54.300 96.300 ;
        RECT 48.500 95.300 50.600 95.600 ;
        RECT 48.500 95.200 48.900 95.300 ;
        RECT 44.600 95.100 45.000 95.200 ;
        RECT 42.500 94.800 45.000 95.100 ;
        RECT 47.000 94.800 47.400 95.200 ;
        RECT 49.300 94.900 49.700 95.000 ;
        RECT 42.500 94.700 42.900 94.800 ;
        RECT 43.800 94.700 44.200 94.800 ;
        RECT 43.300 94.200 43.700 94.300 ;
        RECT 47.000 94.200 47.300 94.800 ;
        RECT 47.800 94.600 49.700 94.900 ;
        RECT 47.800 94.500 48.200 94.600 ;
        RECT 40.600 93.800 41.000 94.200 ;
        RECT 41.800 93.900 47.300 94.200 ;
        RECT 41.800 93.800 42.600 93.900 ;
        RECT 40.600 93.200 40.900 93.800 ;
        RECT 39.800 92.800 40.900 93.200 ;
        RECT 37.400 91.100 37.800 92.200 ;
        RECT 40.300 91.100 40.700 92.800 ;
        RECT 41.400 91.100 41.800 93.500 ;
        RECT 43.900 92.800 44.200 93.900 ;
        RECT 46.700 93.800 47.100 93.900 ;
        RECT 50.200 93.600 50.600 95.300 ;
        RECT 53.500 94.200 53.800 95.900 ;
        RECT 54.200 95.100 54.600 95.600 ;
        RECT 55.000 95.100 55.400 99.900 ;
        RECT 56.600 95.900 57.000 99.900 ;
        RECT 57.400 96.200 57.800 99.900 ;
        RECT 59.000 96.200 59.400 99.900 ;
        RECT 60.600 97.900 61.000 99.900 ;
        RECT 60.700 97.800 61.000 97.900 ;
        RECT 62.200 97.900 62.600 99.900 ;
        RECT 62.200 97.800 62.500 97.900 ;
        RECT 60.700 97.500 62.500 97.800 ;
        RECT 60.600 97.100 61.000 97.200 ;
        RECT 61.400 97.100 61.800 97.200 ;
        RECT 60.600 96.800 61.800 97.100 ;
        RECT 61.400 96.400 61.800 96.800 ;
        RECT 62.200 96.200 62.500 97.500 ;
        RECT 64.300 96.300 64.700 99.900 ;
        RECT 57.400 95.900 59.400 96.200 ;
        RECT 56.700 95.200 57.000 95.900 ;
        RECT 59.800 95.400 60.200 96.200 ;
        RECT 62.200 95.800 62.600 96.200 ;
        RECT 63.800 95.900 64.700 96.300 ;
        RECT 66.700 99.200 67.700 99.900 ;
        RECT 66.700 98.800 68.200 99.200 ;
        RECT 66.700 95.900 67.700 98.800 ;
        RECT 70.700 96.200 71.100 99.900 ;
        RECT 71.400 96.800 71.800 97.200 ;
        RECT 71.500 96.200 71.800 96.800 ;
        RECT 73.900 96.200 74.300 99.900 ;
        RECT 74.600 96.800 75.000 97.200 ;
        RECT 74.700 96.200 75.000 96.800 ;
        RECT 70.700 95.900 71.200 96.200 ;
        RECT 71.500 95.900 72.200 96.200 ;
        RECT 73.900 95.900 74.400 96.200 ;
        RECT 74.700 96.100 75.400 96.200 ;
        RECT 75.800 96.100 76.200 99.900 ;
        RECT 78.500 97.200 78.900 99.900 ;
        RECT 77.800 96.800 78.200 97.200 ;
        RECT 78.500 96.800 79.400 97.200 ;
        RECT 77.800 96.200 78.100 96.800 ;
        RECT 78.500 96.200 78.900 96.800 ;
        RECT 74.700 95.900 76.200 96.100 ;
        RECT 58.600 95.200 59.000 95.400 ;
        RECT 54.200 94.800 55.400 95.100 ;
        RECT 56.600 94.900 57.800 95.200 ;
        RECT 58.600 94.900 59.400 95.200 ;
        RECT 56.600 94.800 57.000 94.900 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 48.700 93.300 50.600 93.600 ;
        RECT 48.700 93.200 49.100 93.300 ;
        RECT 43.000 92.100 43.400 92.500 ;
        RECT 43.800 92.400 44.200 92.800 ;
        RECT 44.700 92.700 45.100 92.800 ;
        RECT 44.700 92.400 46.100 92.700 ;
        RECT 45.800 92.100 46.100 92.400 ;
        RECT 47.800 92.100 48.200 92.500 ;
        RECT 43.000 91.800 44.000 92.100 ;
        RECT 43.600 91.100 44.000 91.800 ;
        RECT 45.800 91.100 46.200 92.100 ;
        RECT 47.800 91.800 48.500 92.100 ;
        RECT 47.900 91.100 48.500 91.800 ;
        RECT 50.200 91.100 50.600 93.300 ;
        RECT 52.600 92.400 53.000 93.200 ;
        RECT 53.500 92.100 53.800 93.800 ;
        RECT 53.400 91.100 53.800 92.100 ;
        RECT 55.000 91.100 55.400 94.800 ;
        RECT 55.800 92.400 56.200 93.200 ;
        RECT 56.600 92.800 57.000 93.200 ;
        RECT 57.500 93.100 57.800 94.900 ;
        RECT 59.000 94.800 59.400 94.900 ;
        RECT 60.600 94.800 61.400 95.200 ;
        RECT 58.200 93.800 58.600 94.600 ;
        RECT 62.200 94.200 62.500 95.800 ;
        RECT 63.900 94.200 64.200 95.900 ;
        RECT 64.600 95.100 65.000 95.600 ;
        RECT 66.200 95.100 66.600 95.200 ;
        RECT 64.600 94.800 66.600 95.100 ;
        RECT 66.200 94.400 66.600 94.800 ;
        RECT 67.000 94.200 67.300 95.900 ;
        RECT 67.800 94.400 68.200 95.200 ;
        RECT 61.700 94.100 62.500 94.200 ;
        RECT 61.600 93.900 62.500 94.100 ;
        RECT 63.000 94.100 63.400 94.200 ;
        RECT 63.800 94.100 64.200 94.200 ;
        RECT 56.700 92.400 57.100 92.800 ;
        RECT 57.400 91.100 57.800 93.100 ;
        RECT 61.600 92.200 62.000 93.900 ;
        RECT 63.000 93.800 64.200 94.100 ;
        RECT 64.600 94.100 65.000 94.200 ;
        RECT 65.400 94.100 65.800 94.200 ;
        RECT 67.000 94.100 67.400 94.200 ;
        RECT 64.600 93.800 66.200 94.100 ;
        RECT 67.000 93.800 68.200 94.100 ;
        RECT 68.600 93.800 69.000 94.600 ;
        RECT 70.200 94.400 70.600 95.200 ;
        RECT 70.900 94.200 71.200 95.900 ;
        RECT 71.800 95.800 72.200 95.900 ;
        RECT 72.600 94.800 73.000 95.200 ;
        RECT 72.600 94.200 72.900 94.800 ;
        RECT 73.400 94.400 73.800 95.200 ;
        RECT 74.100 94.200 74.400 95.900 ;
        RECT 75.000 95.800 76.200 95.900 ;
        RECT 76.600 96.100 77.000 96.200 ;
        RECT 77.400 96.100 78.100 96.200 ;
        RECT 76.600 95.900 78.100 96.100 ;
        RECT 78.400 95.900 78.900 96.200 ;
        RECT 81.900 96.200 82.300 99.900 ;
        RECT 82.600 96.800 83.000 97.200 ;
        RECT 82.700 96.200 83.000 96.800 ;
        RECT 81.900 95.900 82.400 96.200 ;
        RECT 82.700 95.900 83.400 96.200 ;
        RECT 76.600 95.800 77.800 95.900 ;
        RECT 75.000 94.800 75.400 95.200 ;
        RECT 75.000 94.200 75.300 94.800 ;
        RECT 69.400 94.100 69.800 94.200 ;
        RECT 69.400 93.800 70.200 94.100 ;
        RECT 70.900 93.800 72.200 94.200 ;
        RECT 72.600 94.100 73.000 94.200 ;
        RECT 72.600 93.800 73.400 94.100 ;
        RECT 74.100 93.800 75.400 94.200 ;
        RECT 63.000 92.400 63.400 93.200 ;
        RECT 61.400 91.800 62.000 92.200 ;
        RECT 63.900 92.100 64.200 93.800 ;
        RECT 65.800 93.600 66.200 93.800 ;
        RECT 65.500 93.100 67.300 93.300 ;
        RECT 67.900 93.100 68.200 93.800 ;
        RECT 69.800 93.600 70.200 93.800 ;
        RECT 69.500 93.100 71.300 93.300 ;
        RECT 71.800 93.100 72.100 93.800 ;
        RECT 73.000 93.600 73.400 93.800 ;
        RECT 72.700 93.100 74.500 93.300 ;
        RECT 75.000 93.100 75.300 93.800 ;
        RECT 61.600 91.100 62.000 91.800 ;
        RECT 63.800 91.100 64.200 92.100 ;
        RECT 65.400 93.000 67.400 93.100 ;
        RECT 65.400 91.100 65.800 93.000 ;
        RECT 67.000 91.400 67.400 93.000 ;
        RECT 67.800 91.700 68.200 93.100 ;
        RECT 68.600 91.400 69.000 93.100 ;
        RECT 67.000 91.100 69.000 91.400 ;
        RECT 69.400 93.000 71.400 93.100 ;
        RECT 69.400 91.100 69.800 93.000 ;
        RECT 71.000 91.100 71.400 93.000 ;
        RECT 71.800 91.100 72.200 93.100 ;
        RECT 72.600 93.000 74.600 93.100 ;
        RECT 72.600 91.100 73.000 93.000 ;
        RECT 74.200 91.100 74.600 93.000 ;
        RECT 75.000 91.100 75.400 93.100 ;
        RECT 75.800 91.100 76.200 95.800 ;
        RECT 78.400 94.200 78.700 95.900 ;
        RECT 79.000 95.100 79.400 95.200 ;
        RECT 79.800 95.100 80.200 95.200 ;
        RECT 81.400 95.100 81.800 95.200 ;
        RECT 79.000 94.800 81.800 95.100 ;
        RECT 79.000 94.400 79.400 94.800 ;
        RECT 81.400 94.400 81.800 94.800 ;
        RECT 82.100 95.100 82.400 95.900 ;
        RECT 83.000 95.800 83.400 95.900 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 82.100 94.800 83.400 95.100 ;
        RECT 82.100 94.200 82.400 94.800 ;
        RECT 77.400 93.800 78.700 94.200 ;
        RECT 79.800 94.100 80.200 94.200 ;
        RECT 80.600 94.100 81.000 94.200 ;
        RECT 79.400 93.800 81.400 94.100 ;
        RECT 82.100 93.800 83.400 94.200 ;
        RECT 76.600 92.400 77.000 93.200 ;
        RECT 77.500 93.100 77.800 93.800 ;
        RECT 79.400 93.600 79.800 93.800 ;
        RECT 81.000 93.600 81.400 93.800 ;
        RECT 78.300 93.100 80.100 93.300 ;
        RECT 80.700 93.100 82.500 93.300 ;
        RECT 83.000 93.100 83.300 93.800 ;
        RECT 83.800 93.400 84.200 94.200 ;
        RECT 84.600 93.100 85.000 99.900 ;
        RECT 85.400 95.800 85.800 96.600 ;
        RECT 86.200 93.400 86.600 94.200 ;
        RECT 87.000 93.100 87.400 99.900 ;
        RECT 87.800 95.800 88.200 96.600 ;
        RECT 88.600 95.800 89.000 96.600 ;
        RECT 89.400 93.100 89.800 99.900 ;
        RECT 91.800 97.900 92.200 99.900 ;
        RECT 91.900 97.800 92.200 97.900 ;
        RECT 93.400 97.900 93.800 99.900 ;
        RECT 93.400 97.800 93.700 97.900 ;
        RECT 91.900 97.500 93.700 97.800 ;
        RECT 92.600 96.400 93.000 97.200 ;
        RECT 93.400 96.200 93.700 97.500 ;
        RECT 95.000 97.100 95.400 99.900 ;
        RECT 94.200 96.800 95.400 97.100 ;
        RECT 94.200 96.200 94.500 96.800 ;
        RECT 91.000 95.100 91.400 96.200 ;
        RECT 93.400 95.800 93.800 96.200 ;
        RECT 94.200 95.800 94.600 96.200 ;
        RECT 90.200 94.800 91.400 95.100 ;
        RECT 91.800 94.800 92.600 95.200 ;
        RECT 90.200 94.200 90.500 94.800 ;
        RECT 93.400 94.200 93.700 95.800 ;
        RECT 90.200 93.400 90.600 94.200 ;
        RECT 92.900 94.100 93.700 94.200 ;
        RECT 92.800 93.900 93.700 94.100 ;
        RECT 77.400 91.100 77.800 93.100 ;
        RECT 78.200 93.000 80.200 93.100 ;
        RECT 78.200 91.100 78.600 93.000 ;
        RECT 79.800 91.100 80.200 93.000 ;
        RECT 80.600 93.000 82.600 93.100 ;
        RECT 80.600 91.100 81.000 93.000 ;
        RECT 82.200 91.100 82.600 93.000 ;
        RECT 83.000 91.100 83.400 93.100 ;
        RECT 84.600 92.800 85.500 93.100 ;
        RECT 87.000 92.800 87.900 93.100 ;
        RECT 85.100 91.100 85.500 92.800 ;
        RECT 87.500 91.100 87.900 92.800 ;
        RECT 88.900 92.800 89.800 93.100 ;
        RECT 88.900 91.100 89.300 92.800 ;
        RECT 92.800 91.100 93.200 93.900 ;
        RECT 94.200 93.400 94.600 94.200 ;
        RECT 95.000 93.100 95.400 96.800 ;
        RECT 95.800 95.800 96.200 96.600 ;
        RECT 96.600 93.400 97.000 94.200 ;
        RECT 97.400 93.100 97.800 99.900 ;
        RECT 101.900 99.200 102.900 99.900 ;
        RECT 101.400 98.800 102.900 99.200 ;
        RECT 98.200 96.100 98.600 96.600 ;
        RECT 99.000 96.100 99.400 96.200 ;
        RECT 98.200 95.800 99.400 96.100 ;
        RECT 101.900 95.900 102.900 98.800 ;
        RECT 104.600 96.200 105.000 99.900 ;
        RECT 106.200 99.600 108.200 99.900 ;
        RECT 106.200 96.200 106.600 99.600 ;
        RECT 104.600 95.900 106.600 96.200 ;
        RECT 107.000 95.900 107.400 99.300 ;
        RECT 107.800 95.900 108.200 99.600 ;
        RECT 108.600 97.100 109.000 97.200 ;
        RECT 109.400 97.100 109.800 99.900 ;
        RECT 111.800 97.900 112.200 99.900 ;
        RECT 111.900 97.800 112.200 97.900 ;
        RECT 113.400 97.900 113.800 99.900 ;
        RECT 113.400 97.800 113.700 97.900 ;
        RECT 111.900 97.500 113.700 97.800 ;
        RECT 108.600 96.800 109.800 97.100 ;
        RECT 101.400 94.400 101.800 95.200 ;
        RECT 102.200 94.200 102.500 95.900 ;
        RECT 107.000 95.600 107.300 95.900 ;
        RECT 105.000 95.200 105.400 95.400 ;
        RECT 106.300 95.300 107.300 95.600 ;
        RECT 106.300 95.200 106.600 95.300 ;
        RECT 103.000 94.400 103.400 95.200 ;
        RECT 104.600 94.900 105.400 95.200 ;
        RECT 104.600 94.800 105.000 94.900 ;
        RECT 106.200 94.800 106.600 95.200 ;
        RECT 107.800 94.800 108.200 95.600 ;
        RECT 100.600 94.100 101.000 94.200 ;
        RECT 102.200 94.100 102.600 94.200 ;
        RECT 100.600 93.800 101.400 94.100 ;
        RECT 102.200 93.800 103.400 94.100 ;
        RECT 103.800 93.800 104.200 94.600 ;
        RECT 105.400 93.800 105.800 94.600 ;
        RECT 101.000 93.600 101.400 93.800 ;
        RECT 100.700 93.100 102.500 93.300 ;
        RECT 103.100 93.100 103.400 93.800 ;
        RECT 106.300 93.200 106.600 94.800 ;
        RECT 106.900 94.400 107.300 94.800 ;
        RECT 107.000 94.200 107.300 94.400 ;
        RECT 107.000 93.800 107.400 94.200 ;
        RECT 107.800 94.100 108.100 94.800 ;
        RECT 108.600 94.100 109.000 94.200 ;
        RECT 107.800 93.800 109.000 94.100 ;
        RECT 108.600 93.400 109.000 93.800 ;
        RECT 106.200 93.100 106.600 93.200 ;
        RECT 109.400 93.100 109.800 96.800 ;
        RECT 110.200 95.800 110.600 96.600 ;
        RECT 112.600 96.400 113.000 97.200 ;
        RECT 113.400 96.200 113.700 97.500 ;
        RECT 114.200 96.200 114.600 99.900 ;
        RECT 115.800 96.200 116.200 99.900 ;
        RECT 111.000 95.400 111.400 96.200 ;
        RECT 113.400 95.800 113.800 96.200 ;
        RECT 114.200 95.900 116.200 96.200 ;
        RECT 116.600 95.900 117.000 99.900 ;
        RECT 117.700 96.300 118.100 99.900 ;
        RECT 117.700 95.900 118.600 96.300 ;
        RECT 121.100 96.200 121.500 99.900 ;
        RECT 123.800 97.900 124.200 99.900 ;
        RECT 123.900 97.800 124.200 97.900 ;
        RECT 125.400 97.900 125.800 99.900 ;
        RECT 126.200 97.900 126.600 99.900 ;
        RECT 125.400 97.800 125.700 97.900 ;
        RECT 123.900 97.500 125.700 97.800 ;
        RECT 121.800 96.800 122.200 97.200 ;
        RECT 123.800 97.100 124.200 97.200 ;
        RECT 124.600 97.100 125.000 97.200 ;
        RECT 123.800 96.800 125.000 97.100 ;
        RECT 121.900 96.200 122.200 96.800 ;
        RECT 124.600 96.400 125.000 96.800 ;
        RECT 125.400 96.200 125.700 97.500 ;
        RECT 126.300 97.800 126.600 97.900 ;
        RECT 127.800 97.900 128.200 99.900 ;
        RECT 129.400 97.900 129.800 99.900 ;
        RECT 127.800 97.800 128.100 97.900 ;
        RECT 126.300 97.500 128.100 97.800 ;
        RECT 129.500 97.800 129.800 97.900 ;
        RECT 131.000 97.900 131.400 99.900 ;
        RECT 132.600 97.900 133.000 99.900 ;
        RECT 131.000 97.800 131.300 97.900 ;
        RECT 129.500 97.500 131.300 97.800 ;
        RECT 132.700 97.800 133.000 97.900 ;
        RECT 134.200 97.900 134.600 99.900 ;
        RECT 136.600 97.900 137.000 99.900 ;
        RECT 134.200 97.800 134.500 97.900 ;
        RECT 132.700 97.500 134.500 97.800 ;
        RECT 136.700 97.800 137.000 97.900 ;
        RECT 138.200 97.900 138.600 99.900 ;
        RECT 139.800 97.900 140.200 99.900 ;
        RECT 138.200 97.800 138.500 97.900 ;
        RECT 136.700 97.500 138.500 97.800 ;
        RECT 139.900 97.800 140.200 97.900 ;
        RECT 141.400 97.900 141.800 99.900 ;
        RECT 141.400 97.800 141.700 97.900 ;
        RECT 139.900 97.500 141.700 97.800 ;
        RECT 126.300 96.200 126.600 97.500 ;
        RECT 127.000 96.400 127.400 97.200 ;
        RECT 129.500 96.200 129.800 97.500 ;
        RECT 130.200 96.400 130.600 97.200 ;
        RECT 132.700 96.200 133.000 97.500 ;
        RECT 133.400 96.400 133.800 97.200 ;
        RECT 137.400 96.400 137.800 97.200 ;
        RECT 138.200 96.200 138.500 97.500 ;
        RECT 140.600 96.400 141.000 97.200 ;
        RECT 141.400 96.200 141.700 97.500 ;
        RECT 142.200 96.200 142.600 99.900 ;
        RECT 143.800 96.200 144.200 99.900 ;
        RECT 121.100 95.900 121.600 96.200 ;
        RECT 121.900 95.900 122.600 96.200 ;
        RECT 111.800 94.800 112.600 95.200 ;
        RECT 113.400 94.200 113.700 95.800 ;
        RECT 114.600 95.200 115.000 95.400 ;
        RECT 116.600 95.200 116.900 95.900 ;
        RECT 114.200 94.900 115.000 95.200 ;
        RECT 115.800 94.900 117.000 95.200 ;
        RECT 114.200 94.800 114.600 94.900 ;
        RECT 115.800 94.800 116.200 94.900 ;
        RECT 116.600 94.800 117.000 94.900 ;
        RECT 117.400 94.800 117.800 95.600 ;
        RECT 112.900 94.100 113.700 94.200 ;
        RECT 112.800 93.900 113.700 94.100 ;
        RECT 95.000 92.800 95.900 93.100 ;
        RECT 97.400 92.800 98.300 93.100 ;
        RECT 95.500 91.100 95.900 92.800 ;
        RECT 97.900 91.100 98.300 92.800 ;
        RECT 100.600 93.000 102.600 93.100 ;
        RECT 100.600 91.100 101.000 93.000 ;
        RECT 102.200 91.400 102.600 93.000 ;
        RECT 103.000 91.700 103.400 93.100 ;
        RECT 103.800 91.400 104.200 93.100 ;
        RECT 102.200 91.100 104.200 91.400 ;
        RECT 106.100 91.100 106.900 93.100 ;
        RECT 109.400 92.800 110.300 93.100 ;
        RECT 109.900 91.100 110.300 92.800 ;
        RECT 112.800 91.100 113.200 93.900 ;
        RECT 115.000 93.800 115.400 94.600 ;
        RECT 115.800 93.100 116.100 94.800 ;
        RECT 118.200 94.200 118.500 95.900 ;
        RECT 119.800 95.100 120.200 95.200 ;
        RECT 120.600 95.100 121.000 95.200 ;
        RECT 119.800 94.800 121.000 95.100 ;
        RECT 120.600 94.400 121.000 94.800 ;
        RECT 121.300 95.100 121.600 95.900 ;
        RECT 122.200 95.800 122.600 95.900 ;
        RECT 123.000 95.400 123.400 96.200 ;
        RECT 125.400 95.800 125.800 96.200 ;
        RECT 126.200 95.800 126.600 96.200 ;
        RECT 122.200 95.100 122.600 95.200 ;
        RECT 121.300 94.800 122.600 95.100 ;
        RECT 123.800 94.800 124.600 95.200 ;
        RECT 121.300 94.200 121.600 94.800 ;
        RECT 125.400 94.200 125.700 95.800 ;
        RECT 118.200 94.100 118.600 94.200 ;
        RECT 119.800 94.100 120.200 94.200 ;
        RECT 118.200 93.800 120.600 94.100 ;
        RECT 121.300 93.800 122.600 94.200 ;
        RECT 124.900 94.100 125.700 94.200 ;
        RECT 124.800 93.900 125.700 94.100 ;
        RECT 126.300 94.200 126.600 95.800 ;
        RECT 128.600 95.400 129.000 96.200 ;
        RECT 129.400 95.800 129.800 96.200 ;
        RECT 127.400 94.800 128.200 95.200 ;
        RECT 129.500 94.200 129.800 95.800 ;
        RECT 131.800 95.400 132.200 96.200 ;
        RECT 132.600 95.800 133.000 96.200 ;
        RECT 134.200 96.100 134.600 96.200 ;
        RECT 135.000 96.100 135.400 96.200 ;
        RECT 135.800 96.100 136.200 96.200 ;
        RECT 134.200 95.800 136.200 96.100 ;
        RECT 130.600 94.800 131.400 95.200 ;
        RECT 132.700 94.200 133.000 95.800 ;
        RECT 135.000 95.400 135.400 95.800 ;
        RECT 135.800 95.400 136.200 95.800 ;
        RECT 138.200 95.800 138.600 96.200 ;
        RECT 133.800 94.800 134.600 95.200 ;
        RECT 136.600 94.800 137.400 95.200 ;
        RECT 138.200 94.200 138.500 95.800 ;
        RECT 139.000 95.400 139.400 96.200 ;
        RECT 141.400 95.800 141.800 96.200 ;
        RECT 142.200 95.900 144.200 96.200 ;
        RECT 144.600 95.900 145.000 99.900 ;
        RECT 139.800 94.800 140.600 95.200 ;
        RECT 141.400 95.100 141.700 95.800 ;
        RECT 142.600 95.200 143.000 95.400 ;
        RECT 144.600 95.200 144.900 95.900 ;
        RECT 142.200 95.100 143.000 95.200 ;
        RECT 141.400 94.900 143.000 95.100 ;
        RECT 143.800 94.900 145.000 95.200 ;
        RECT 141.400 94.800 142.600 94.900 ;
        RECT 141.400 94.200 141.700 94.800 ;
        RECT 126.300 94.100 127.100 94.200 ;
        RECT 129.500 94.100 130.300 94.200 ;
        RECT 132.700 94.100 133.500 94.200 ;
        RECT 137.700 94.100 138.500 94.200 ;
        RECT 140.900 94.100 141.700 94.200 ;
        RECT 126.300 93.900 127.200 94.100 ;
        RECT 129.500 93.900 130.400 94.100 ;
        RECT 132.700 93.900 134.500 94.100 ;
        RECT 115.800 91.100 116.200 93.100 ;
        RECT 116.600 92.800 117.000 93.200 ;
        RECT 116.500 92.400 116.900 92.800 ;
        RECT 118.200 92.100 118.500 93.800 ;
        RECT 120.200 93.600 120.600 93.800 ;
        RECT 119.000 92.400 119.400 93.200 ;
        RECT 119.900 93.100 121.700 93.300 ;
        RECT 122.200 93.100 122.500 93.800 ;
        RECT 119.800 93.000 121.800 93.100 ;
        RECT 118.200 91.100 118.600 92.100 ;
        RECT 119.800 91.100 120.200 93.000 ;
        RECT 121.400 91.100 121.800 93.000 ;
        RECT 122.200 91.100 122.600 93.100 ;
        RECT 124.800 91.100 125.200 93.900 ;
        RECT 126.800 91.100 127.200 93.900 ;
        RECT 130.000 92.200 130.400 93.900 ;
        RECT 133.200 93.800 134.500 93.900 ;
        RECT 130.000 91.800 130.600 92.200 ;
        RECT 130.000 91.100 130.400 91.800 ;
        RECT 133.200 91.100 133.600 93.800 ;
        RECT 134.200 93.200 134.500 93.800 ;
        RECT 137.600 93.900 138.500 94.100 ;
        RECT 140.800 93.900 141.700 94.100 ;
        RECT 134.200 92.800 134.600 93.200 ;
        RECT 136.600 92.100 137.000 92.200 ;
        RECT 137.600 92.100 138.000 93.900 ;
        RECT 136.600 91.800 138.000 92.100 ;
        RECT 137.600 91.100 138.000 91.800 ;
        RECT 140.800 92.200 141.200 93.900 ;
        RECT 143.000 93.800 143.400 94.600 ;
        RECT 143.800 93.100 144.100 94.900 ;
        RECT 144.600 94.800 145.000 94.900 ;
        RECT 145.400 93.400 145.800 94.200 ;
        RECT 140.800 91.800 141.800 92.200 ;
        RECT 140.800 91.100 141.200 91.800 ;
        RECT 143.800 91.100 144.200 93.100 ;
        RECT 144.600 92.800 145.000 93.200 ;
        RECT 146.200 93.100 146.600 99.900 ;
        RECT 147.800 97.900 148.200 99.900 ;
        RECT 147.900 97.800 148.200 97.900 ;
        RECT 149.400 97.900 149.800 99.900 ;
        RECT 149.400 97.800 149.700 97.900 ;
        RECT 147.900 97.500 149.700 97.800 ;
        RECT 147.000 95.800 147.400 96.600 ;
        RECT 147.900 96.200 148.200 97.500 ;
        RECT 148.600 96.400 149.000 97.200 ;
        RECT 147.800 95.800 148.200 96.200 ;
        RECT 147.000 94.800 147.400 95.200 ;
        RECT 147.000 94.100 147.300 94.800 ;
        RECT 147.900 94.200 148.200 95.800 ;
        RECT 150.200 95.400 150.600 96.200 ;
        RECT 149.000 94.800 149.800 95.200 ;
        RECT 147.900 94.100 148.700 94.200 ;
        RECT 147.000 93.800 148.800 94.100 ;
        RECT 146.200 92.800 147.100 93.100 ;
        RECT 144.500 92.400 144.900 92.800 ;
        RECT 146.700 92.200 147.100 92.800 ;
        RECT 146.200 91.800 147.100 92.200 ;
        RECT 146.700 91.100 147.100 91.800 ;
        RECT 148.400 91.100 148.800 93.800 ;
        RECT 1.400 85.100 1.800 89.900 ;
        RECT 3.500 88.200 3.900 89.900 ;
        RECT 5.400 88.900 5.800 89.900 ;
        RECT 3.000 87.900 3.900 88.200 ;
        RECT 1.400 84.800 2.500 85.100 ;
        RECT 1.400 81.100 1.800 84.800 ;
        RECT 2.200 84.200 2.500 84.800 ;
        RECT 2.200 83.800 2.600 84.200 ;
        RECT 3.000 81.100 3.400 87.900 ;
        RECT 4.600 87.800 5.000 88.600 ;
        RECT 5.500 87.800 5.800 88.900 ;
        RECT 7.000 87.900 7.400 89.900 ;
        RECT 7.800 87.900 8.200 89.900 ;
        RECT 9.900 89.200 10.300 89.900 ;
        RECT 9.900 88.800 10.600 89.200 ;
        RECT 9.900 88.400 10.300 88.800 ;
        RECT 9.900 87.900 10.600 88.400 ;
        RECT 11.000 87.900 11.400 89.900 ;
        RECT 11.800 88.000 12.200 89.900 ;
        RECT 13.400 88.000 13.800 89.900 ;
        RECT 11.800 87.900 13.800 88.000 ;
        RECT 3.800 87.100 4.200 87.200 ;
        RECT 4.600 87.100 4.900 87.800 ;
        RECT 5.500 87.500 6.700 87.800 ;
        RECT 3.800 86.800 4.900 87.100 ;
        RECT 6.400 86.000 6.700 87.500 ;
        RECT 7.100 87.100 7.400 87.900 ;
        RECT 7.900 87.800 8.200 87.900 ;
        RECT 7.900 87.600 8.800 87.800 ;
        RECT 7.900 87.500 10.000 87.600 ;
        RECT 8.500 87.300 10.000 87.500 ;
        RECT 9.600 87.200 10.000 87.300 ;
        RECT 7.800 87.100 8.200 87.200 ;
        RECT 7.000 86.800 8.200 87.100 ;
        RECT 8.800 86.900 9.200 87.000 ;
        RECT 7.100 86.200 7.400 86.800 ;
        RECT 7.800 86.400 8.200 86.800 ;
        RECT 8.700 86.600 9.200 86.900 ;
        RECT 8.700 86.200 9.000 86.600 ;
        RECT 6.300 85.700 6.700 86.000 ;
        RECT 7.000 85.800 7.400 86.200 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 4.600 85.600 6.700 85.700 ;
        RECT 4.600 85.400 6.600 85.600 ;
        RECT 3.800 84.400 4.200 85.200 ;
        RECT 4.600 81.100 5.000 85.400 ;
        RECT 7.100 85.100 7.400 85.800 ;
        RECT 9.600 85.500 9.900 87.200 ;
        RECT 10.300 86.200 10.600 87.900 ;
        RECT 11.100 87.200 11.400 87.900 ;
        RECT 11.900 87.700 13.700 87.900 ;
        RECT 14.200 87.800 14.600 88.600 ;
        RECT 13.000 87.200 13.400 87.400 ;
        RECT 11.000 86.800 12.300 87.200 ;
        RECT 13.000 87.100 13.800 87.200 ;
        RECT 15.000 87.100 15.400 89.900 ;
        RECT 15.900 88.200 16.300 88.600 ;
        RECT 13.000 86.900 15.400 87.100 ;
        RECT 13.400 86.800 15.400 86.900 ;
        RECT 15.800 87.800 16.200 88.200 ;
        RECT 16.600 87.900 17.000 89.900 ;
        RECT 19.800 88.900 20.200 89.900 ;
        RECT 15.800 87.200 16.100 87.800 ;
        RECT 15.800 86.800 16.200 87.200 ;
        RECT 10.200 85.800 10.600 86.200 ;
        RECT 8.700 85.200 9.900 85.500 ;
        RECT 6.700 84.800 8.100 85.100 ;
        RECT 6.700 81.100 7.100 84.800 ;
        RECT 7.800 84.200 8.100 84.800 ;
        RECT 7.800 83.800 8.200 84.200 ;
        RECT 8.700 83.100 9.000 85.200 ;
        RECT 10.300 85.100 10.600 85.800 ;
        RECT 8.600 81.100 9.000 83.100 ;
        RECT 10.200 81.100 10.600 85.100 ;
        RECT 11.000 85.100 11.400 85.200 ;
        RECT 12.000 85.100 12.300 86.800 ;
        RECT 12.600 85.800 13.000 86.600 ;
        RECT 11.000 84.800 11.700 85.100 ;
        RECT 12.000 84.800 12.500 85.100 ;
        RECT 11.400 84.200 11.700 84.800 ;
        RECT 11.400 83.800 11.800 84.200 ;
        RECT 12.100 82.200 12.500 84.800 ;
        RECT 12.100 81.800 13.000 82.200 ;
        RECT 12.100 81.100 12.500 81.800 ;
        RECT 15.000 81.100 15.400 86.800 ;
        RECT 15.800 86.100 16.200 86.200 ;
        RECT 16.700 86.100 17.000 87.900 ;
        RECT 19.000 87.800 19.400 88.600 ;
        RECT 19.900 87.200 20.200 88.900 ;
        RECT 17.400 86.400 17.800 87.200 ;
        RECT 19.800 86.800 20.200 87.200 ;
        RECT 21.400 86.800 21.800 87.600 ;
        RECT 22.200 87.100 22.600 89.900 ;
        RECT 23.000 87.900 23.400 89.900 ;
        RECT 25.200 89.200 26.000 89.900 ;
        RECT 24.600 88.800 26.000 89.200 ;
        RECT 25.200 88.100 26.000 88.800 ;
        RECT 23.000 87.600 24.200 87.900 ;
        RECT 23.800 87.500 24.200 87.600 ;
        RECT 24.500 87.400 24.900 87.800 ;
        RECT 24.500 87.200 24.800 87.400 ;
        RECT 23.000 87.100 23.800 87.200 ;
        RECT 22.200 86.800 23.800 87.100 ;
        RECT 24.400 86.800 24.800 87.200 ;
        RECT 18.200 86.100 18.600 86.200 ;
        RECT 15.800 85.800 17.000 86.100 ;
        RECT 17.800 85.800 18.600 86.100 ;
        RECT 15.900 85.100 16.200 85.800 ;
        RECT 17.800 85.600 18.200 85.800 ;
        RECT 19.900 85.100 20.200 86.800 ;
        RECT 20.600 86.100 21.000 86.200 ;
        RECT 22.200 86.100 22.600 86.800 ;
        RECT 25.200 86.400 25.500 88.100 ;
        RECT 27.800 87.900 28.200 89.900 ;
        RECT 25.800 87.700 26.600 87.800 ;
        RECT 25.800 87.400 26.800 87.700 ;
        RECT 27.100 87.600 28.200 87.900 ;
        RECT 27.100 87.500 27.500 87.600 ;
        RECT 28.600 87.500 29.000 89.900 ;
        RECT 30.800 89.200 31.200 89.900 ;
        RECT 30.200 88.900 31.200 89.200 ;
        RECT 33.000 88.900 33.400 89.900 ;
        RECT 35.100 89.200 35.700 89.900 ;
        RECT 35.000 88.900 35.700 89.200 ;
        RECT 30.200 88.500 30.600 88.900 ;
        RECT 33.000 88.600 33.300 88.900 ;
        RECT 31.000 87.800 31.400 88.600 ;
        RECT 31.900 88.300 33.300 88.600 ;
        RECT 35.000 88.500 35.400 88.900 ;
        RECT 31.900 88.200 32.300 88.300 ;
        RECT 26.500 87.200 26.800 87.400 ;
        RECT 25.800 86.700 26.200 87.100 ;
        RECT 26.500 86.900 28.200 87.200 ;
        RECT 27.400 86.800 28.200 86.900 ;
        RECT 29.000 87.100 29.800 87.200 ;
        RECT 31.100 87.100 31.400 87.800 ;
        RECT 35.900 87.700 36.300 87.800 ;
        RECT 37.400 87.700 37.800 89.900 ;
        RECT 35.900 87.400 37.800 87.700 ;
        RECT 38.200 87.500 38.600 89.900 ;
        RECT 40.400 89.200 40.800 89.900 ;
        RECT 39.800 88.900 40.800 89.200 ;
        RECT 42.600 88.900 43.000 89.900 ;
        RECT 44.700 89.200 45.300 89.900 ;
        RECT 44.600 88.900 45.300 89.200 ;
        RECT 39.800 88.500 40.200 88.900 ;
        RECT 42.600 88.600 42.900 88.900 ;
        RECT 40.600 88.200 41.000 88.600 ;
        RECT 41.500 88.300 42.900 88.600 ;
        RECT 44.600 88.500 45.000 88.900 ;
        RECT 41.500 88.200 41.900 88.300 ;
        RECT 33.900 87.100 34.300 87.200 ;
        RECT 29.000 86.800 34.500 87.100 ;
        RECT 30.500 86.700 30.900 86.800 ;
        RECT 25.000 86.200 25.500 86.400 ;
        RECT 20.600 85.800 22.600 86.100 ;
        RECT 24.600 86.100 25.500 86.200 ;
        RECT 25.900 86.400 26.200 86.700 ;
        RECT 25.900 86.100 27.200 86.400 ;
        RECT 24.600 85.800 25.300 86.100 ;
        RECT 26.800 86.000 27.200 86.100 ;
        RECT 29.700 86.200 30.100 86.300 ;
        RECT 31.000 86.200 31.400 86.300 ;
        RECT 29.700 85.900 32.200 86.200 ;
        RECT 31.800 85.800 32.200 85.900 ;
        RECT 20.600 85.400 21.000 85.800 ;
        RECT 15.800 81.100 16.200 85.100 ;
        RECT 16.600 84.800 18.600 85.100 ;
        RECT 16.600 81.100 17.000 84.800 ;
        RECT 18.200 81.100 18.600 84.800 ;
        RECT 19.800 84.700 20.700 85.100 ;
        RECT 20.300 82.200 20.700 84.700 ;
        RECT 19.800 81.800 20.700 82.200 ;
        RECT 20.300 81.100 20.700 81.800 ;
        RECT 22.200 81.100 22.600 85.800 ;
        RECT 25.000 85.100 25.300 85.800 ;
        RECT 25.700 85.700 26.100 85.800 ;
        RECT 25.700 85.400 27.400 85.700 ;
        RECT 27.100 85.100 27.400 85.400 ;
        RECT 28.600 85.500 31.400 85.600 ;
        RECT 28.600 85.400 31.500 85.500 ;
        RECT 28.600 85.300 33.500 85.400 ;
        RECT 23.000 84.800 24.200 85.100 ;
        RECT 25.000 84.800 26.000 85.100 ;
        RECT 23.000 81.100 23.400 84.800 ;
        RECT 23.800 84.700 24.200 84.800 ;
        RECT 25.200 81.100 26.000 84.800 ;
        RECT 27.100 84.800 28.200 85.100 ;
        RECT 27.100 84.700 27.500 84.800 ;
        RECT 27.800 81.100 28.200 84.800 ;
        RECT 28.600 81.100 29.000 85.300 ;
        RECT 31.100 85.100 33.500 85.300 ;
        RECT 30.200 84.500 32.900 84.800 ;
        RECT 30.200 84.400 30.600 84.500 ;
        RECT 32.500 84.400 32.900 84.500 ;
        RECT 33.200 84.500 33.500 85.100 ;
        RECT 34.200 85.200 34.500 86.800 ;
        RECT 35.000 86.400 35.400 86.500 ;
        RECT 35.000 86.100 36.900 86.400 ;
        RECT 36.500 86.000 36.900 86.100 ;
        RECT 35.700 85.700 36.100 85.800 ;
        RECT 37.400 85.700 37.800 87.400 ;
        RECT 38.600 87.100 39.400 87.200 ;
        RECT 40.700 87.100 41.000 88.200 ;
        RECT 45.500 87.700 45.900 87.800 ;
        RECT 47.000 87.700 47.400 89.900 ;
        RECT 45.500 87.400 47.400 87.700 ;
        RECT 49.400 87.500 49.800 89.900 ;
        RECT 51.600 89.200 52.000 89.900 ;
        RECT 51.000 88.900 52.000 89.200 ;
        RECT 53.800 88.900 54.200 89.900 ;
        RECT 55.900 89.200 56.500 89.900 ;
        RECT 55.800 88.900 56.500 89.200 ;
        RECT 51.000 88.500 51.400 88.900 ;
        RECT 53.800 88.600 54.100 88.900 ;
        RECT 51.800 88.200 52.200 88.600 ;
        RECT 52.700 88.300 54.100 88.600 ;
        RECT 55.800 88.500 56.200 88.900 ;
        RECT 52.700 88.200 53.100 88.300 ;
        RECT 43.500 87.100 43.900 87.200 ;
        RECT 38.600 86.800 44.100 87.100 ;
        RECT 40.100 86.700 40.500 86.800 ;
        RECT 43.000 86.100 43.400 86.200 ;
        RECT 43.800 86.100 44.100 86.800 ;
        RECT 44.600 86.400 45.000 86.500 ;
        RECT 44.600 86.100 46.500 86.400 ;
        RECT 43.000 85.800 44.100 86.100 ;
        RECT 46.100 86.000 46.500 86.100 ;
        RECT 47.000 86.100 47.400 87.400 ;
        RECT 49.800 87.100 50.600 87.200 ;
        RECT 51.900 87.100 52.200 88.200 ;
        RECT 56.700 87.700 57.100 87.800 ;
        RECT 58.200 87.700 58.600 89.900 ;
        RECT 59.000 87.800 59.400 88.600 ;
        RECT 56.700 87.400 58.600 87.700 ;
        RECT 54.700 87.100 55.100 87.200 ;
        RECT 49.800 86.800 55.300 87.100 ;
        RECT 51.300 86.700 51.700 86.800 ;
        RECT 50.500 86.200 50.900 86.300 ;
        RECT 51.800 86.200 52.200 86.300 ;
        RECT 47.800 86.100 48.200 86.200 ;
        RECT 47.000 85.800 48.200 86.100 ;
        RECT 50.500 85.900 53.000 86.200 ;
        RECT 52.600 85.800 53.000 85.900 ;
        RECT 35.700 85.400 37.800 85.700 ;
        RECT 34.200 84.900 35.400 85.200 ;
        RECT 33.900 84.500 34.300 84.600 ;
        RECT 33.200 84.200 34.300 84.500 ;
        RECT 35.100 84.400 35.400 84.900 ;
        RECT 35.100 84.000 35.800 84.400 ;
        RECT 31.900 83.700 32.300 83.800 ;
        RECT 33.300 83.700 33.700 83.800 ;
        RECT 30.200 83.100 30.600 83.500 ;
        RECT 31.900 83.400 33.700 83.700 ;
        RECT 33.000 83.100 33.300 83.400 ;
        RECT 35.000 83.100 35.400 83.500 ;
        RECT 30.200 82.800 31.200 83.100 ;
        RECT 30.800 81.100 31.200 82.800 ;
        RECT 33.000 81.100 33.400 83.100 ;
        RECT 35.100 81.100 35.700 83.100 ;
        RECT 37.400 81.100 37.800 85.400 ;
        RECT 38.200 85.500 41.000 85.600 ;
        RECT 38.200 85.400 41.100 85.500 ;
        RECT 38.200 85.300 43.100 85.400 ;
        RECT 38.200 81.100 38.600 85.300 ;
        RECT 40.700 85.100 43.100 85.300 ;
        RECT 39.800 84.500 42.500 84.800 ;
        RECT 39.800 84.400 40.200 84.500 ;
        RECT 42.100 84.400 42.500 84.500 ;
        RECT 42.800 84.500 43.100 85.100 ;
        RECT 43.800 85.200 44.100 85.800 ;
        RECT 45.300 85.700 45.700 85.800 ;
        RECT 47.000 85.700 47.400 85.800 ;
        RECT 45.300 85.400 47.400 85.700 ;
        RECT 43.800 84.900 45.000 85.200 ;
        RECT 43.500 84.500 43.900 84.600 ;
        RECT 42.800 84.200 43.900 84.500 ;
        RECT 44.700 84.400 45.000 84.900 ;
        RECT 44.700 84.000 45.400 84.400 ;
        RECT 41.500 83.700 41.900 83.800 ;
        RECT 42.900 83.700 43.300 83.800 ;
        RECT 39.800 83.100 40.200 83.500 ;
        RECT 41.500 83.400 43.300 83.700 ;
        RECT 42.600 83.100 42.900 83.400 ;
        RECT 44.600 83.100 45.000 83.500 ;
        RECT 39.800 82.800 40.800 83.100 ;
        RECT 40.400 81.100 40.800 82.800 ;
        RECT 42.600 81.100 43.000 83.100 ;
        RECT 44.700 81.100 45.300 83.100 ;
        RECT 47.000 81.100 47.400 85.400 ;
        RECT 49.400 85.500 52.200 85.600 ;
        RECT 49.400 85.400 52.300 85.500 ;
        RECT 49.400 85.300 54.300 85.400 ;
        RECT 49.400 81.100 49.800 85.300 ;
        RECT 51.900 85.100 54.300 85.300 ;
        RECT 51.000 84.500 53.700 84.800 ;
        RECT 51.000 84.400 51.400 84.500 ;
        RECT 53.300 84.400 53.700 84.500 ;
        RECT 54.000 84.500 54.300 85.100 ;
        RECT 55.000 85.200 55.300 86.800 ;
        RECT 55.800 86.400 56.200 86.500 ;
        RECT 55.800 86.100 57.700 86.400 ;
        RECT 57.300 86.000 57.700 86.100 ;
        RECT 56.500 85.700 56.900 85.800 ;
        RECT 58.200 85.700 58.600 87.400 ;
        RECT 56.500 85.400 58.600 85.700 ;
        RECT 55.000 84.900 56.200 85.200 ;
        RECT 54.700 84.500 55.100 84.600 ;
        RECT 54.000 84.200 55.100 84.500 ;
        RECT 55.900 84.400 56.200 84.900 ;
        RECT 55.900 84.000 56.600 84.400 ;
        RECT 52.700 83.700 53.100 83.800 ;
        RECT 54.100 83.700 54.500 83.800 ;
        RECT 51.000 83.100 51.400 83.500 ;
        RECT 52.700 83.400 54.500 83.700 ;
        RECT 53.800 83.100 54.100 83.400 ;
        RECT 55.800 83.100 56.200 83.500 ;
        RECT 51.000 82.800 52.000 83.100 ;
        RECT 51.600 81.100 52.000 82.800 ;
        RECT 53.800 81.100 54.200 83.100 ;
        RECT 55.900 81.100 56.500 83.100 ;
        RECT 58.200 81.100 58.600 85.400 ;
        RECT 59.800 87.100 60.200 89.900 ;
        RECT 60.600 87.900 61.000 89.900 ;
        RECT 62.700 89.200 63.100 89.900 ;
        RECT 65.100 89.200 65.500 89.900 ;
        RECT 67.500 89.200 67.900 89.900 ;
        RECT 68.900 89.200 69.300 89.900 ;
        RECT 62.700 88.800 63.400 89.200 ;
        RECT 65.100 88.800 65.800 89.200 ;
        RECT 67.000 88.800 67.900 89.200 ;
        RECT 68.600 88.800 69.300 89.200 ;
        RECT 62.700 88.400 63.100 88.800 ;
        RECT 62.700 87.900 63.400 88.400 ;
        RECT 65.100 88.200 65.500 88.800 ;
        RECT 67.500 88.200 67.900 88.800 ;
        RECT 60.700 87.800 61.000 87.900 ;
        RECT 60.700 87.600 61.600 87.800 ;
        RECT 60.700 87.500 62.800 87.600 ;
        RECT 61.300 87.300 62.800 87.500 ;
        RECT 62.400 87.200 62.800 87.300 ;
        RECT 60.600 87.100 61.000 87.200 ;
        RECT 59.800 86.800 61.000 87.100 ;
        RECT 61.600 86.900 62.000 87.000 ;
        RECT 59.800 81.100 60.200 86.800 ;
        RECT 60.600 86.400 61.000 86.800 ;
        RECT 61.500 86.600 62.000 86.900 ;
        RECT 61.500 86.200 61.800 86.600 ;
        RECT 61.400 85.800 61.800 86.200 ;
        RECT 62.400 85.500 62.700 87.200 ;
        RECT 63.100 86.200 63.400 87.900 ;
        RECT 64.600 87.900 65.500 88.200 ;
        RECT 67.000 87.900 67.900 88.200 ;
        RECT 68.900 88.200 69.300 88.800 ;
        RECT 68.900 87.900 69.800 88.200 ;
        RECT 72.300 87.900 73.100 89.900 ;
        RECT 76.300 89.200 76.700 89.900 ;
        RECT 76.300 88.800 77.000 89.200 ;
        RECT 76.300 88.200 76.700 88.800 ;
        RECT 78.700 88.200 79.100 89.900 ;
        RECT 79.900 88.200 80.300 88.600 ;
        RECT 75.800 87.900 76.700 88.200 ;
        RECT 78.200 88.100 79.100 88.200 ;
        RECT 79.800 88.100 80.200 88.200 ;
        RECT 63.800 86.800 64.200 87.600 ;
        RECT 63.000 85.800 63.400 86.200 ;
        RECT 61.500 85.200 62.700 85.500 ;
        RECT 61.500 83.100 61.800 85.200 ;
        RECT 63.100 85.100 63.400 85.800 ;
        RECT 61.400 81.100 61.800 83.100 ;
        RECT 63.000 81.100 63.400 85.100 ;
        RECT 64.600 81.100 65.000 87.900 ;
        RECT 66.200 86.800 66.600 87.600 ;
        RECT 65.400 85.100 65.800 85.200 ;
        RECT 66.200 85.100 66.600 85.200 ;
        RECT 65.400 84.800 66.600 85.100 ;
        RECT 65.400 84.400 65.800 84.800 ;
        RECT 67.000 81.100 67.400 87.900 ;
        RECT 67.800 84.400 68.200 85.200 ;
        RECT 68.600 84.400 69.000 85.200 ;
        RECT 69.400 81.100 69.800 87.900 ;
        RECT 70.200 87.100 70.600 87.600 ;
        RECT 70.200 86.800 71.300 87.100 ;
        RECT 71.800 86.800 72.200 87.200 ;
        RECT 71.000 86.200 71.300 86.800 ;
        RECT 71.900 86.600 72.200 86.800 ;
        RECT 71.900 86.200 72.300 86.600 ;
        RECT 72.600 86.200 72.900 87.900 ;
        RECT 73.400 86.400 73.800 87.200 ;
        RECT 75.000 87.100 75.400 87.600 ;
        RECT 74.200 86.800 75.400 87.100 ;
        RECT 74.200 86.200 74.500 86.800 ;
        RECT 71.000 85.400 71.400 86.200 ;
        RECT 72.600 85.800 73.000 86.200 ;
        RECT 74.200 86.100 74.600 86.200 ;
        RECT 73.800 85.800 74.600 86.100 ;
        RECT 72.600 85.700 72.900 85.800 ;
        RECT 71.900 85.400 72.900 85.700 ;
        RECT 73.800 85.600 74.200 85.800 ;
        RECT 71.900 85.100 72.200 85.400 ;
        RECT 71.000 81.400 71.400 85.100 ;
        RECT 71.800 81.700 72.200 85.100 ;
        RECT 72.600 84.800 74.600 85.100 ;
        RECT 72.600 81.400 73.000 84.800 ;
        RECT 71.000 81.100 73.000 81.400 ;
        RECT 74.200 81.100 74.600 84.800 ;
        RECT 75.800 81.100 76.200 87.900 ;
        RECT 78.200 87.800 80.200 88.100 ;
        RECT 80.600 87.900 81.000 89.900 ;
        RECT 77.400 86.800 77.800 87.600 ;
        RECT 76.600 84.400 77.000 85.200 ;
        RECT 78.200 81.100 78.600 87.800 ;
        RECT 79.800 86.100 80.200 86.200 ;
        RECT 80.700 86.100 81.000 87.900 ;
        RECT 81.400 86.400 81.800 87.200 ;
        RECT 82.200 87.100 82.600 87.200 ;
        RECT 83.000 87.100 83.400 89.900 ;
        RECT 83.800 87.800 84.200 88.600 ;
        RECT 86.200 87.900 86.600 89.900 ;
        RECT 86.900 88.200 87.300 88.600 ;
        RECT 89.100 88.200 89.500 89.900 ;
        RECT 82.200 86.800 83.400 87.100 ;
        RECT 83.800 87.100 84.200 87.200 ;
        RECT 85.400 87.100 85.800 87.200 ;
        RECT 83.800 86.800 85.800 87.100 ;
        RECT 82.200 86.100 82.600 86.200 ;
        RECT 79.800 85.800 81.000 86.100 ;
        RECT 81.800 85.800 82.600 86.100 ;
        RECT 79.000 84.400 79.400 85.200 ;
        RECT 79.900 85.100 80.200 85.800 ;
        RECT 81.800 85.600 82.200 85.800 ;
        RECT 79.800 81.100 80.200 85.100 ;
        RECT 80.600 84.800 82.600 85.100 ;
        RECT 80.600 81.100 81.000 84.800 ;
        RECT 82.200 81.100 82.600 84.800 ;
        RECT 83.000 81.100 83.400 86.800 ;
        RECT 85.400 86.400 85.800 86.800 ;
        RECT 84.600 86.100 85.000 86.200 ;
        RECT 86.200 86.100 86.500 87.900 ;
        RECT 87.000 87.800 87.400 88.200 ;
        RECT 88.600 87.900 89.500 88.200 ;
        RECT 87.000 87.100 87.400 87.200 ;
        RECT 87.800 87.100 88.200 87.600 ;
        RECT 87.000 86.800 88.200 87.100 ;
        RECT 87.000 86.100 87.400 86.200 ;
        RECT 84.600 85.800 85.400 86.100 ;
        RECT 86.200 85.800 87.400 86.100 ;
        RECT 85.000 85.600 85.400 85.800 ;
        RECT 87.000 85.100 87.300 85.800 ;
        RECT 84.600 84.800 86.600 85.100 ;
        RECT 84.600 81.100 85.000 84.800 ;
        RECT 86.200 81.100 86.600 84.800 ;
        RECT 87.000 81.100 87.400 85.100 ;
        RECT 88.600 81.100 89.000 87.900 ;
        RECT 90.200 87.800 90.600 88.600 ;
        RECT 91.000 86.100 91.400 89.900 ;
        RECT 91.800 88.000 92.200 89.900 ;
        RECT 93.400 88.000 93.800 89.900 ;
        RECT 91.800 87.900 93.800 88.000 ;
        RECT 94.200 87.900 94.600 89.900 ;
        RECT 96.300 87.900 97.100 89.900 ;
        RECT 100.300 88.200 100.700 89.900 ;
        RECT 103.300 89.200 103.700 89.900 ;
        RECT 103.000 88.800 103.700 89.200 ;
        RECT 99.800 87.900 100.700 88.200 ;
        RECT 103.300 88.200 103.700 88.800 ;
        RECT 103.300 87.900 104.200 88.200 ;
        RECT 91.900 87.700 93.700 87.900 ;
        RECT 92.200 87.200 92.600 87.400 ;
        RECT 94.200 87.200 94.500 87.900 ;
        RECT 91.800 86.900 92.600 87.200 ;
        RECT 93.300 87.100 94.600 87.200 ;
        RECT 95.000 87.100 95.400 87.200 ;
        RECT 91.800 86.800 92.200 86.900 ;
        RECT 93.300 86.800 95.400 87.100 ;
        RECT 95.800 86.800 96.200 87.200 ;
        RECT 92.600 86.100 93.000 86.600 ;
        RECT 91.000 85.800 93.000 86.100 ;
        RECT 89.400 84.400 89.800 85.200 ;
        RECT 91.000 81.100 91.400 85.800 ;
        RECT 93.300 85.100 93.600 86.800 ;
        RECT 95.900 86.600 96.200 86.800 ;
        RECT 95.900 86.200 96.300 86.600 ;
        RECT 96.600 86.200 96.900 87.900 ;
        RECT 97.400 86.400 97.800 87.200 ;
        RECT 99.000 86.800 99.400 87.600 ;
        RECT 95.000 85.400 95.400 86.200 ;
        RECT 96.600 85.800 97.000 86.200 ;
        RECT 98.200 86.100 98.600 86.200 ;
        RECT 97.800 85.800 98.600 86.100 ;
        RECT 96.600 85.700 96.900 85.800 ;
        RECT 95.900 85.400 96.900 85.700 ;
        RECT 97.800 85.600 98.200 85.800 ;
        RECT 94.200 85.100 94.600 85.200 ;
        RECT 95.900 85.100 96.200 85.400 ;
        RECT 93.100 84.800 93.600 85.100 ;
        RECT 93.900 84.800 94.600 85.100 ;
        RECT 93.100 81.100 93.500 84.800 ;
        RECT 93.900 84.200 94.200 84.800 ;
        RECT 93.800 83.800 94.200 84.200 ;
        RECT 95.000 81.400 95.400 85.100 ;
        RECT 95.800 81.700 96.200 85.100 ;
        RECT 96.600 84.800 98.600 85.100 ;
        RECT 96.600 81.400 97.000 84.800 ;
        RECT 95.000 81.100 97.000 81.400 ;
        RECT 98.200 81.100 98.600 84.800 ;
        RECT 99.800 81.100 100.200 87.900 ;
        RECT 100.600 84.400 101.000 85.200 ;
        RECT 101.400 85.100 101.800 85.200 ;
        RECT 103.000 85.100 103.400 85.200 ;
        RECT 101.400 84.800 103.400 85.100 ;
        RECT 103.000 84.400 103.400 84.800 ;
        RECT 103.800 84.100 104.200 87.900 ;
        RECT 104.600 86.800 105.000 87.600 ;
        RECT 107.200 87.100 107.600 89.900 ;
        RECT 110.200 87.900 110.600 89.900 ;
        RECT 110.900 88.200 111.300 88.600 ;
        RECT 107.200 86.900 108.100 87.100 ;
        RECT 107.300 86.800 108.100 86.900 ;
        RECT 106.200 85.800 107.000 86.200 ;
        RECT 105.400 84.800 105.800 85.600 ;
        RECT 107.800 85.200 108.100 86.800 ;
        RECT 109.400 86.400 109.800 87.200 ;
        RECT 108.600 86.100 109.000 86.200 ;
        RECT 110.200 86.100 110.500 87.900 ;
        RECT 111.000 87.800 111.400 88.200 ;
        RECT 111.000 86.800 111.400 87.200 ;
        RECT 113.600 87.100 114.000 89.900 ;
        RECT 116.600 87.900 117.000 89.900 ;
        RECT 117.300 88.200 117.700 88.600 ;
        RECT 116.600 87.200 116.900 87.900 ;
        RECT 117.400 87.800 117.800 88.200 ;
        RECT 118.200 88.000 118.600 89.900 ;
        RECT 119.800 89.600 121.800 89.900 ;
        RECT 119.800 88.000 120.200 89.600 ;
        RECT 118.200 87.900 120.200 88.000 ;
        RECT 120.600 87.900 121.000 89.300 ;
        RECT 121.400 87.900 121.800 89.600 ;
        RECT 123.000 88.900 123.400 89.900 ;
        RECT 118.300 87.700 120.100 87.900 ;
        RECT 118.600 87.200 119.000 87.400 ;
        RECT 120.700 87.200 121.000 87.900 ;
        RECT 122.200 87.800 122.600 88.600 ;
        RECT 123.100 87.200 123.400 88.900 ;
        RECT 124.600 87.900 125.000 89.900 ;
        RECT 125.400 88.000 125.800 89.900 ;
        RECT 127.000 88.000 127.400 89.900 ;
        RECT 125.400 87.900 127.400 88.000 ;
        RECT 127.800 88.000 128.200 89.900 ;
        RECT 129.400 88.000 129.800 89.900 ;
        RECT 127.800 87.900 129.800 88.000 ;
        RECT 130.200 87.900 130.600 89.900 ;
        RECT 131.100 88.200 131.500 88.600 ;
        RECT 124.700 87.200 125.000 87.900 ;
        RECT 125.500 87.700 127.300 87.900 ;
        RECT 127.900 87.700 129.700 87.900 ;
        RECT 126.600 87.200 127.000 87.400 ;
        RECT 128.200 87.200 128.600 87.400 ;
        RECT 130.200 87.200 130.500 87.900 ;
        RECT 131.000 87.800 131.400 88.200 ;
        RECT 131.800 87.900 132.200 89.900 ;
        RECT 113.600 86.900 114.500 87.100 ;
        RECT 113.700 86.800 114.500 86.900 ;
        RECT 111.000 86.200 111.300 86.800 ;
        RECT 111.000 86.100 111.400 86.200 ;
        RECT 108.600 85.800 109.400 86.100 ;
        RECT 110.200 85.800 111.400 86.100 ;
        RECT 112.600 85.800 113.400 86.200 ;
        RECT 109.000 85.600 109.400 85.800 ;
        RECT 107.000 84.100 107.400 85.200 ;
        RECT 103.800 83.800 107.400 84.100 ;
        RECT 107.800 84.800 108.200 85.200 ;
        RECT 111.000 85.100 111.300 85.800 ;
        RECT 108.600 84.800 110.600 85.100 ;
        RECT 103.800 81.100 104.200 83.800 ;
        RECT 107.800 83.500 108.100 84.800 ;
        RECT 106.300 83.200 108.100 83.500 ;
        RECT 106.300 83.100 106.600 83.200 ;
        RECT 106.200 81.100 106.600 83.100 ;
        RECT 107.800 83.100 108.100 83.200 ;
        RECT 107.800 81.100 108.200 83.100 ;
        RECT 108.600 81.100 109.000 84.800 ;
        RECT 110.200 81.100 110.600 84.800 ;
        RECT 111.000 81.100 111.400 85.100 ;
        RECT 111.800 84.800 112.200 85.600 ;
        RECT 114.200 85.200 114.500 86.800 ;
        RECT 115.800 86.400 116.200 87.200 ;
        RECT 116.600 86.800 117.000 87.200 ;
        RECT 118.200 86.900 119.000 87.200 ;
        RECT 119.800 86.900 121.000 87.200 ;
        RECT 118.200 86.800 118.600 86.900 ;
        RECT 119.800 86.800 120.200 86.900 ;
        RECT 115.000 86.100 115.400 86.200 ;
        RECT 116.600 86.100 116.900 86.800 ;
        RECT 117.400 86.100 117.800 86.200 ;
        RECT 115.000 85.800 115.800 86.100 ;
        RECT 116.600 85.800 117.800 86.100 ;
        RECT 119.000 85.800 119.400 86.600 ;
        RECT 115.400 85.600 115.800 85.800 ;
        RECT 114.200 84.800 114.600 85.200 ;
        RECT 117.400 85.100 117.700 85.800 ;
        RECT 119.800 85.100 120.100 86.800 ;
        RECT 120.600 85.800 121.000 86.600 ;
        RECT 121.400 86.400 121.800 87.200 ;
        RECT 123.000 86.800 123.400 87.200 ;
        RECT 124.600 86.800 125.900 87.200 ;
        RECT 126.600 87.100 127.400 87.200 ;
        RECT 127.800 87.100 128.600 87.200 ;
        RECT 126.600 86.900 128.600 87.100 ;
        RECT 127.000 86.800 128.200 86.900 ;
        RECT 129.300 86.800 130.600 87.200 ;
        RECT 123.100 85.100 123.400 86.800 ;
        RECT 123.800 85.400 124.200 86.200 ;
        RECT 124.600 85.100 125.000 85.200 ;
        RECT 125.600 85.100 125.900 86.800 ;
        RECT 126.200 86.100 126.600 86.600 ;
        RECT 128.600 86.100 129.000 86.600 ;
        RECT 126.200 85.800 129.000 86.100 ;
        RECT 129.300 85.100 129.600 86.800 ;
        RECT 131.000 86.100 131.400 86.200 ;
        RECT 131.900 86.100 132.200 87.900 ;
        RECT 132.600 86.400 133.000 87.200 ;
        RECT 134.800 87.100 135.200 89.900 ;
        RECT 138.000 87.100 138.400 89.900 ;
        RECT 142.200 87.900 142.600 89.900 ;
        RECT 142.900 88.200 143.300 88.600 ;
        RECT 134.300 86.900 135.200 87.100 ;
        RECT 137.500 86.900 138.400 87.100 ;
        RECT 134.300 86.800 135.100 86.900 ;
        RECT 137.500 86.800 138.300 86.900 ;
        RECT 133.400 86.100 133.800 86.200 ;
        RECT 131.000 85.800 132.200 86.100 ;
        RECT 133.000 85.800 133.800 86.100 ;
        RECT 130.200 85.100 130.600 85.200 ;
        RECT 131.100 85.100 131.400 85.800 ;
        RECT 133.000 85.600 133.400 85.800 ;
        RECT 134.300 85.200 134.600 86.800 ;
        RECT 135.400 85.800 136.200 86.200 ;
        RECT 115.000 84.800 117.000 85.100 ;
        RECT 113.400 83.800 113.800 84.600 ;
        RECT 114.200 83.500 114.500 84.800 ;
        RECT 112.700 83.200 114.500 83.500 ;
        RECT 112.700 83.100 113.000 83.200 ;
        RECT 112.600 81.100 113.000 83.100 ;
        RECT 114.200 83.100 114.500 83.200 ;
        RECT 114.200 81.100 114.600 83.100 ;
        RECT 115.000 81.100 115.400 84.800 ;
        RECT 116.600 81.100 117.000 84.800 ;
        RECT 117.400 81.100 117.800 85.100 ;
        RECT 119.500 81.100 120.500 85.100 ;
        RECT 123.000 84.700 123.900 85.100 ;
        RECT 124.600 84.800 125.300 85.100 ;
        RECT 125.600 84.800 126.100 85.100 ;
        RECT 123.500 84.200 123.900 84.700 ;
        RECT 125.000 84.200 125.300 84.800 ;
        RECT 123.500 83.800 124.200 84.200 ;
        RECT 125.000 83.800 125.400 84.200 ;
        RECT 123.500 81.100 123.900 83.800 ;
        RECT 125.700 82.200 126.100 84.800 ;
        RECT 129.100 84.800 129.600 85.100 ;
        RECT 129.900 84.800 130.600 85.100 ;
        RECT 129.100 82.200 129.500 84.800 ;
        RECT 129.900 84.200 130.200 84.800 ;
        RECT 129.800 83.800 130.200 84.200 ;
        RECT 125.700 81.800 126.600 82.200 ;
        RECT 128.600 81.800 129.500 82.200 ;
        RECT 125.700 81.100 126.100 81.800 ;
        RECT 129.100 81.100 129.500 81.800 ;
        RECT 131.000 81.100 131.400 85.100 ;
        RECT 131.800 84.800 133.800 85.100 ;
        RECT 134.200 84.800 134.600 85.200 ;
        RECT 136.600 84.800 137.000 85.600 ;
        RECT 137.500 85.200 137.800 86.800 ;
        RECT 141.400 86.400 141.800 87.200 ;
        RECT 138.600 85.800 139.400 86.200 ;
        RECT 140.600 86.100 141.000 86.200 ;
        RECT 142.200 86.100 142.500 87.900 ;
        RECT 143.000 87.800 143.400 88.200 ;
        RECT 145.600 87.100 146.000 89.900 ;
        RECT 148.800 87.100 149.200 89.900 ;
        RECT 145.600 86.900 146.500 87.100 ;
        RECT 148.800 86.900 149.700 87.100 ;
        RECT 145.700 86.800 146.500 86.900 ;
        RECT 148.900 86.800 149.700 86.900 ;
        RECT 143.000 86.100 143.400 86.200 ;
        RECT 139.800 85.800 141.400 86.100 ;
        RECT 142.200 85.800 143.400 86.100 ;
        RECT 144.600 85.800 145.400 86.200 ;
        RECT 137.400 84.800 137.800 85.200 ;
        RECT 139.800 84.800 140.200 85.800 ;
        RECT 141.000 85.600 141.400 85.800 ;
        RECT 143.000 85.100 143.300 85.800 ;
        RECT 140.600 84.800 142.600 85.100 ;
        RECT 131.800 81.100 132.200 84.800 ;
        RECT 133.400 81.100 133.800 84.800 ;
        RECT 134.300 83.500 134.600 84.800 ;
        RECT 135.000 83.800 135.400 84.600 ;
        RECT 137.500 83.500 137.800 84.800 ;
        RECT 138.200 83.800 138.600 84.600 ;
        RECT 134.300 83.200 136.100 83.500 ;
        RECT 134.300 83.100 134.600 83.200 ;
        RECT 134.200 81.100 134.600 83.100 ;
        RECT 135.800 83.100 136.100 83.200 ;
        RECT 137.500 83.200 139.300 83.500 ;
        RECT 137.500 83.100 137.800 83.200 ;
        RECT 135.800 81.100 136.200 83.100 ;
        RECT 137.400 81.100 137.800 83.100 ;
        RECT 139.000 83.100 139.300 83.200 ;
        RECT 139.000 81.100 139.400 83.100 ;
        RECT 140.600 81.100 141.000 84.800 ;
        RECT 142.200 81.100 142.600 84.800 ;
        RECT 143.000 81.100 143.400 85.100 ;
        RECT 143.800 84.800 144.200 85.600 ;
        RECT 146.200 85.200 146.500 86.800 ;
        RECT 147.800 85.800 148.600 86.200 ;
        RECT 146.200 84.800 146.600 85.200 ;
        RECT 147.000 84.800 147.400 85.600 ;
        RECT 149.400 85.200 149.700 86.800 ;
        RECT 149.400 84.800 149.800 85.200 ;
        RECT 145.400 83.800 145.800 84.600 ;
        RECT 146.200 83.500 146.500 84.800 ;
        RECT 148.600 83.800 149.000 84.600 ;
        RECT 149.400 83.500 149.700 84.800 ;
        RECT 144.700 83.200 146.500 83.500 ;
        RECT 144.700 83.100 145.000 83.200 ;
        RECT 144.600 81.100 145.000 83.100 ;
        RECT 146.200 83.100 146.500 83.200 ;
        RECT 147.900 83.200 149.700 83.500 ;
        RECT 147.900 83.100 148.200 83.200 ;
        RECT 146.200 81.100 146.600 83.100 ;
        RECT 147.800 81.100 148.200 83.100 ;
        RECT 149.400 83.100 149.700 83.200 ;
        RECT 149.400 81.100 149.800 83.100 ;
        RECT 1.400 71.100 1.800 79.900 ;
        RECT 3.000 75.100 3.400 79.900 ;
        RECT 5.100 76.300 5.500 79.900 ;
        RECT 4.600 75.900 5.500 76.300 ;
        RECT 6.200 76.200 6.600 79.900 ;
        RECT 6.900 76.200 7.300 76.300 ;
        RECT 6.200 75.900 7.300 76.200 ;
        RECT 8.400 76.200 9.200 79.900 ;
        RECT 10.200 76.200 10.600 76.300 ;
        RECT 11.000 76.200 11.400 79.900 ;
        RECT 8.400 75.900 9.400 76.200 ;
        RECT 10.200 75.900 11.400 76.200 ;
        RECT 3.000 74.800 4.100 75.100 ;
        RECT 3.000 71.100 3.400 74.800 ;
        RECT 3.800 74.200 4.100 74.800 ;
        RECT 4.700 74.200 5.000 75.900 ;
        RECT 7.000 75.600 7.300 75.900 ;
        RECT 5.400 74.800 5.800 75.600 ;
        RECT 7.000 75.300 8.700 75.600 ;
        RECT 8.300 75.200 8.700 75.300 ;
        RECT 9.100 75.200 9.400 75.900 ;
        RECT 7.200 74.900 7.600 75.000 ;
        RECT 9.100 74.900 9.800 75.200 ;
        RECT 7.200 74.600 8.500 74.900 ;
        RECT 3.800 73.800 4.200 74.200 ;
        RECT 4.600 73.800 5.000 74.200 ;
        RECT 8.200 74.300 8.500 74.600 ;
        RECT 8.900 74.800 9.800 74.900 ;
        RECT 8.900 74.600 9.400 74.800 ;
        RECT 8.200 73.900 8.600 74.300 ;
        RECT 3.800 72.400 4.200 73.200 ;
        RECT 4.700 72.200 5.000 73.800 ;
        RECT 6.900 73.400 7.300 73.500 ;
        RECT 4.600 71.100 5.000 72.200 ;
        RECT 6.200 73.100 7.300 73.400 ;
        RECT 6.200 71.100 6.600 73.100 ;
        RECT 8.900 72.900 9.200 74.600 ;
        RECT 12.600 74.100 13.000 79.900 ;
        RECT 14.700 76.200 15.100 79.900 ;
        RECT 15.400 76.800 15.800 77.200 ;
        RECT 15.500 76.200 15.800 76.800 ;
        RECT 14.700 75.900 15.200 76.200 ;
        RECT 15.500 75.900 16.200 76.200 ;
        RECT 16.600 75.900 17.000 79.900 ;
        RECT 17.400 76.200 17.800 79.900 ;
        RECT 19.000 76.200 19.400 79.900 ;
        RECT 17.400 75.900 19.400 76.200 ;
        RECT 14.900 75.200 15.200 75.900 ;
        RECT 15.800 75.800 16.200 75.900 ;
        RECT 16.700 75.200 17.000 75.900 ;
        RECT 19.800 75.700 20.200 79.900 ;
        RECT 22.000 78.200 22.400 79.900 ;
        RECT 21.400 77.900 22.400 78.200 ;
        RECT 24.200 77.900 24.600 79.900 ;
        RECT 26.300 77.900 26.900 79.900 ;
        RECT 21.400 77.500 21.800 77.900 ;
        RECT 24.200 77.600 24.500 77.900 ;
        RECT 23.100 77.300 24.900 77.600 ;
        RECT 26.200 77.500 26.600 77.900 ;
        RECT 23.100 77.200 23.500 77.300 ;
        RECT 24.500 77.200 24.900 77.300 ;
        RECT 21.400 76.500 21.800 76.600 ;
        RECT 23.700 76.500 24.100 76.600 ;
        RECT 21.400 76.200 24.100 76.500 ;
        RECT 24.400 76.500 25.500 76.800 ;
        RECT 24.400 75.900 24.700 76.500 ;
        RECT 25.100 76.400 25.500 76.500 ;
        RECT 26.300 76.600 27.000 77.000 ;
        RECT 26.300 76.100 26.600 76.600 ;
        RECT 22.300 75.700 24.700 75.900 ;
        RECT 19.800 75.600 24.700 75.700 ;
        RECT 25.400 75.800 26.600 76.100 ;
        RECT 19.800 75.500 22.700 75.600 ;
        RECT 19.800 75.400 22.600 75.500 ;
        RECT 18.600 75.200 19.000 75.400 ;
        RECT 14.900 74.800 15.400 75.200 ;
        RECT 16.600 74.900 17.800 75.200 ;
        RECT 18.600 74.900 19.400 75.200 ;
        RECT 16.600 74.800 17.000 74.900 ;
        RECT 14.900 74.200 15.200 74.800 ;
        RECT 13.400 74.100 13.800 74.200 ;
        RECT 12.600 73.800 14.200 74.100 ;
        RECT 14.900 73.800 16.200 74.200 ;
        RECT 10.200 73.400 10.600 73.500 ;
        RECT 10.200 73.100 11.400 73.400 ;
        RECT 8.400 72.200 9.200 72.900 ;
        RECT 8.400 71.800 9.800 72.200 ;
        RECT 8.400 71.100 9.200 71.800 ;
        RECT 11.000 71.100 11.400 73.100 ;
        RECT 12.600 71.100 13.000 73.800 ;
        RECT 13.800 73.600 14.200 73.800 ;
        RECT 13.500 73.100 15.300 73.300 ;
        RECT 15.800 73.100 16.100 73.800 ;
        RECT 13.400 73.000 15.400 73.100 ;
        RECT 13.400 71.100 13.800 73.000 ;
        RECT 15.000 71.100 15.400 73.000 ;
        RECT 15.800 71.100 16.200 73.100 ;
        RECT 16.600 72.800 17.000 73.200 ;
        RECT 17.500 73.100 17.800 74.900 ;
        RECT 19.000 74.800 19.400 74.900 ;
        RECT 18.200 73.800 18.600 74.600 ;
        RECT 21.700 74.200 22.100 74.300 ;
        RECT 25.400 74.200 25.700 75.800 ;
        RECT 28.600 75.600 29.000 79.900 ;
        RECT 26.900 75.300 29.000 75.600 ;
        RECT 29.400 75.700 29.800 79.900 ;
        RECT 31.600 78.200 32.000 79.900 ;
        RECT 31.000 77.900 32.000 78.200 ;
        RECT 33.800 77.900 34.200 79.900 ;
        RECT 35.900 77.900 36.500 79.900 ;
        RECT 31.000 77.500 31.400 77.900 ;
        RECT 33.800 77.600 34.100 77.900 ;
        RECT 32.700 77.300 34.500 77.600 ;
        RECT 35.800 77.500 36.200 77.900 ;
        RECT 32.700 77.200 33.100 77.300 ;
        RECT 34.100 77.200 34.500 77.300 ;
        RECT 31.000 76.500 31.400 76.600 ;
        RECT 33.300 76.500 33.700 76.600 ;
        RECT 31.000 76.200 33.700 76.500 ;
        RECT 34.000 76.500 35.100 76.800 ;
        RECT 34.000 75.900 34.300 76.500 ;
        RECT 34.700 76.400 35.100 76.500 ;
        RECT 35.900 76.600 36.600 77.000 ;
        RECT 35.900 76.100 36.200 76.600 ;
        RECT 31.900 75.700 34.300 75.900 ;
        RECT 29.400 75.600 34.300 75.700 ;
        RECT 35.000 75.800 36.200 76.100 ;
        RECT 29.400 75.500 32.300 75.600 ;
        RECT 29.400 75.400 32.200 75.500 ;
        RECT 26.900 75.200 27.300 75.300 ;
        RECT 27.700 74.900 28.100 75.000 ;
        RECT 26.200 74.600 28.100 74.900 ;
        RECT 26.200 74.500 26.600 74.600 ;
        RECT 20.200 73.900 25.700 74.200 ;
        RECT 20.200 73.800 21.000 73.900 ;
        RECT 16.700 72.400 17.100 72.800 ;
        RECT 17.400 71.100 17.800 73.100 ;
        RECT 19.800 71.100 20.200 73.500 ;
        RECT 22.300 72.800 22.600 73.900 ;
        RECT 25.100 73.800 25.500 73.900 ;
        RECT 28.600 73.600 29.000 75.300 ;
        RECT 35.000 75.200 35.300 75.800 ;
        RECT 38.200 75.600 38.600 79.900 ;
        RECT 36.500 75.300 38.600 75.600 ;
        RECT 39.000 75.700 39.400 79.900 ;
        RECT 41.200 78.200 41.600 79.900 ;
        RECT 40.600 77.900 41.600 78.200 ;
        RECT 43.400 77.900 43.800 79.900 ;
        RECT 45.500 77.900 46.100 79.900 ;
        RECT 40.600 77.500 41.000 77.900 ;
        RECT 43.400 77.600 43.700 77.900 ;
        RECT 42.300 77.300 44.100 77.600 ;
        RECT 45.400 77.500 45.800 77.900 ;
        RECT 42.300 77.200 42.700 77.300 ;
        RECT 43.700 77.200 44.100 77.300 ;
        RECT 40.600 76.500 41.000 76.600 ;
        RECT 42.900 76.500 43.300 76.600 ;
        RECT 40.600 76.200 43.300 76.500 ;
        RECT 43.600 76.500 44.700 76.800 ;
        RECT 43.600 75.900 43.900 76.500 ;
        RECT 44.300 76.400 44.700 76.500 ;
        RECT 45.500 76.600 46.200 77.000 ;
        RECT 45.500 76.100 45.800 76.600 ;
        RECT 41.500 75.700 43.900 75.900 ;
        RECT 39.000 75.600 43.900 75.700 ;
        RECT 44.600 75.800 45.800 76.100 ;
        RECT 39.000 75.500 41.900 75.600 ;
        RECT 39.000 75.400 41.800 75.500 ;
        RECT 36.500 75.200 36.900 75.300 ;
        RECT 35.000 74.800 35.400 75.200 ;
        RECT 37.300 74.900 37.700 75.000 ;
        RECT 31.300 74.200 31.700 74.300 ;
        RECT 35.000 74.200 35.300 74.800 ;
        RECT 35.800 74.600 37.700 74.900 ;
        RECT 35.800 74.500 36.200 74.600 ;
        RECT 29.800 73.900 35.300 74.200 ;
        RECT 29.800 73.800 30.600 73.900 ;
        RECT 27.100 73.300 29.000 73.600 ;
        RECT 27.100 73.200 27.500 73.300 ;
        RECT 21.400 72.100 21.800 72.500 ;
        RECT 22.200 72.400 22.600 72.800 ;
        RECT 23.100 72.700 23.500 72.800 ;
        RECT 23.100 72.400 24.500 72.700 ;
        RECT 24.200 72.100 24.500 72.400 ;
        RECT 26.200 72.100 26.600 72.500 ;
        RECT 21.400 71.800 22.400 72.100 ;
        RECT 22.000 71.100 22.400 71.800 ;
        RECT 24.200 71.100 24.600 72.100 ;
        RECT 26.200 71.800 26.900 72.100 ;
        RECT 26.300 71.100 26.900 71.800 ;
        RECT 28.600 71.100 29.000 73.300 ;
        RECT 29.400 71.100 29.800 73.500 ;
        RECT 31.900 72.800 32.200 73.900 ;
        RECT 34.700 73.800 35.100 73.900 ;
        RECT 38.200 73.600 38.600 75.300 ;
        RECT 42.200 75.100 42.600 75.200 ;
        RECT 40.100 74.800 42.600 75.100 ;
        RECT 40.100 74.700 40.500 74.800 ;
        RECT 41.400 74.700 41.800 74.800 ;
        RECT 40.900 74.200 41.300 74.300 ;
        RECT 44.600 74.200 44.900 75.800 ;
        RECT 47.800 75.600 48.200 79.900 ;
        RECT 46.100 75.300 48.200 75.600 ;
        RECT 50.200 75.700 50.600 79.900 ;
        RECT 52.400 78.200 52.800 79.900 ;
        RECT 51.800 77.900 52.800 78.200 ;
        RECT 54.600 77.900 55.000 79.900 ;
        RECT 56.700 77.900 57.300 79.900 ;
        RECT 51.800 77.500 52.200 77.900 ;
        RECT 54.600 77.600 54.900 77.900 ;
        RECT 53.500 77.300 55.300 77.600 ;
        RECT 56.600 77.500 57.000 77.900 ;
        RECT 53.500 77.200 53.900 77.300 ;
        RECT 54.900 77.200 55.300 77.300 ;
        RECT 51.800 76.500 52.200 76.600 ;
        RECT 54.100 76.500 54.500 76.600 ;
        RECT 51.800 76.200 54.500 76.500 ;
        RECT 54.800 76.500 55.900 76.800 ;
        RECT 54.800 75.900 55.100 76.500 ;
        RECT 55.500 76.400 55.900 76.500 ;
        RECT 56.700 76.600 57.400 77.000 ;
        RECT 56.700 76.100 57.000 76.600 ;
        RECT 52.700 75.700 55.100 75.900 ;
        RECT 50.200 75.600 55.100 75.700 ;
        RECT 55.800 75.800 57.000 76.100 ;
        RECT 50.200 75.500 53.100 75.600 ;
        RECT 50.200 75.400 53.000 75.500 ;
        RECT 46.100 75.200 46.500 75.300 ;
        RECT 46.900 74.900 47.300 75.000 ;
        RECT 45.400 74.600 47.300 74.900 ;
        RECT 45.400 74.500 45.800 74.600 ;
        RECT 39.400 73.900 44.900 74.200 ;
        RECT 39.400 73.800 40.200 73.900 ;
        RECT 36.700 73.300 38.600 73.600 ;
        RECT 36.700 73.200 37.100 73.300 ;
        RECT 31.000 72.100 31.400 72.500 ;
        RECT 31.800 72.400 32.200 72.800 ;
        RECT 32.700 72.700 33.100 72.800 ;
        RECT 32.700 72.400 34.100 72.700 ;
        RECT 33.800 72.100 34.100 72.400 ;
        RECT 35.800 72.100 36.200 72.500 ;
        RECT 31.000 71.800 32.000 72.100 ;
        RECT 31.600 71.100 32.000 71.800 ;
        RECT 33.800 71.100 34.200 72.100 ;
        RECT 35.800 71.800 36.500 72.100 ;
        RECT 35.900 71.100 36.500 71.800 ;
        RECT 38.200 71.100 38.600 73.300 ;
        RECT 39.000 71.100 39.400 73.500 ;
        RECT 41.500 72.800 41.800 73.900 ;
        RECT 43.000 73.800 43.400 73.900 ;
        RECT 44.300 73.800 44.700 73.900 ;
        RECT 47.800 73.600 48.200 75.300 ;
        RECT 53.400 75.100 53.800 75.200 ;
        RECT 51.300 74.800 53.800 75.100 ;
        RECT 51.300 74.700 51.700 74.800 ;
        RECT 52.600 74.700 53.000 74.800 ;
        RECT 52.100 74.200 52.500 74.300 ;
        RECT 55.800 74.200 56.100 75.800 ;
        RECT 59.000 75.600 59.400 79.900 ;
        RECT 59.800 77.100 60.200 77.200 ;
        RECT 60.600 77.100 61.000 79.900 ;
        RECT 62.200 77.900 62.600 79.900 ;
        RECT 59.800 76.800 61.000 77.100 ;
        RECT 57.300 75.300 59.400 75.600 ;
        RECT 57.300 75.200 57.700 75.300 ;
        RECT 58.100 74.900 58.500 75.000 ;
        RECT 56.600 74.600 58.500 74.900 ;
        RECT 56.600 74.500 57.000 74.600 ;
        RECT 50.600 73.900 56.100 74.200 ;
        RECT 50.600 73.800 51.400 73.900 ;
        RECT 46.300 73.300 48.200 73.600 ;
        RECT 46.300 73.200 46.700 73.300 ;
        RECT 40.600 72.100 41.000 72.500 ;
        RECT 41.400 72.400 41.800 72.800 ;
        RECT 42.300 72.700 42.700 72.800 ;
        RECT 42.300 72.400 43.700 72.700 ;
        RECT 43.400 72.100 43.700 72.400 ;
        RECT 45.400 72.100 45.800 72.500 ;
        RECT 40.600 71.800 41.600 72.100 ;
        RECT 41.200 71.100 41.600 71.800 ;
        RECT 43.400 71.100 43.800 72.100 ;
        RECT 45.400 71.800 46.100 72.100 ;
        RECT 45.500 71.100 46.100 71.800 ;
        RECT 47.800 71.100 48.200 73.300 ;
        RECT 50.200 71.100 50.600 73.500 ;
        RECT 52.700 73.200 53.000 73.900 ;
        RECT 55.500 73.800 55.900 73.900 ;
        RECT 59.000 73.600 59.400 75.300 ;
        RECT 57.500 73.300 59.400 73.600 ;
        RECT 59.800 73.400 60.200 74.200 ;
        RECT 57.500 73.200 57.900 73.300 ;
        RECT 51.800 72.100 52.200 72.500 ;
        RECT 52.600 72.400 53.000 73.200 ;
        RECT 53.500 72.700 53.900 72.800 ;
        RECT 53.500 72.400 54.900 72.700 ;
        RECT 54.600 72.100 54.900 72.400 ;
        RECT 56.600 72.100 57.000 72.500 ;
        RECT 51.800 71.800 52.800 72.100 ;
        RECT 52.400 71.100 52.800 71.800 ;
        RECT 54.600 71.100 55.000 72.100 ;
        RECT 56.600 71.800 57.300 72.100 ;
        RECT 56.700 71.100 57.300 71.800 ;
        RECT 59.000 71.100 59.400 73.300 ;
        RECT 60.600 73.100 61.000 76.800 ;
        RECT 62.300 77.800 62.600 77.900 ;
        RECT 63.800 77.800 64.200 79.900 ;
        RECT 62.300 77.500 64.100 77.800 ;
        RECT 61.400 75.800 61.800 76.600 ;
        RECT 62.300 76.200 62.600 77.500 ;
        RECT 63.000 77.100 63.400 77.200 ;
        RECT 64.600 77.100 65.000 77.200 ;
        RECT 63.000 76.800 65.000 77.100 ;
        RECT 63.000 76.400 63.400 76.800 ;
        RECT 62.200 75.800 62.600 76.200 ;
        RECT 62.300 74.200 62.600 75.800 ;
        RECT 64.600 75.400 65.000 76.200 ;
        RECT 65.400 75.900 65.800 79.900 ;
        RECT 66.200 76.200 66.600 79.900 ;
        RECT 67.800 76.200 68.200 79.900 ;
        RECT 66.200 75.900 68.200 76.200 ;
        RECT 65.500 75.200 65.800 75.900 ;
        RECT 67.400 75.200 67.800 75.400 ;
        RECT 63.400 74.800 64.200 75.200 ;
        RECT 65.400 74.900 66.600 75.200 ;
        RECT 67.400 74.900 68.200 75.200 ;
        RECT 65.400 74.800 65.800 74.900 ;
        RECT 62.300 74.100 63.100 74.200 ;
        RECT 62.300 73.900 63.200 74.100 ;
        RECT 60.600 72.800 61.500 73.100 ;
        RECT 61.100 71.100 61.500 72.800 ;
        RECT 62.800 71.100 63.200 73.900 ;
        RECT 65.400 72.800 65.800 73.200 ;
        RECT 66.300 73.100 66.600 74.900 ;
        RECT 67.800 74.800 68.200 74.900 ;
        RECT 67.000 73.800 67.400 74.600 ;
        RECT 67.800 74.100 68.100 74.800 ;
        RECT 68.600 74.100 69.000 74.200 ;
        RECT 67.800 73.800 69.000 74.100 ;
        RECT 68.600 73.400 69.000 73.800 ;
        RECT 65.500 72.400 65.900 72.800 ;
        RECT 66.200 71.100 66.600 73.100 ;
        RECT 69.400 73.100 69.800 79.900 ;
        RECT 70.200 75.800 70.600 76.600 ;
        RECT 71.000 75.900 71.400 79.900 ;
        RECT 71.800 76.200 72.200 79.900 ;
        RECT 73.400 76.200 73.800 79.900 ;
        RECT 71.800 75.900 73.800 76.200 ;
        RECT 74.200 76.200 74.600 79.900 ;
        RECT 75.800 76.400 76.200 79.900 ;
        RECT 74.200 75.900 75.500 76.200 ;
        RECT 75.800 75.900 76.300 76.400 ;
        RECT 77.400 76.200 77.800 79.900 ;
        RECT 79.000 76.400 79.400 79.900 ;
        RECT 77.400 75.900 78.700 76.200 ;
        RECT 79.000 75.900 79.500 76.400 ;
        RECT 80.600 76.200 81.000 79.900 ;
        RECT 82.200 76.400 82.600 79.900 ;
        RECT 80.600 75.900 81.900 76.200 ;
        RECT 82.200 75.900 82.700 76.400 ;
        RECT 71.100 75.200 71.400 75.900 ;
        RECT 73.000 75.200 73.400 75.400 ;
        RECT 71.000 74.900 72.200 75.200 ;
        RECT 73.000 74.900 73.800 75.200 ;
        RECT 71.000 74.800 71.400 74.900 ;
        RECT 71.800 74.800 72.200 74.900 ;
        RECT 73.400 74.800 73.800 74.900 ;
        RECT 74.200 74.800 74.700 75.200 ;
        RECT 71.000 73.100 71.400 73.200 ;
        RECT 71.900 73.100 72.200 74.800 ;
        RECT 72.600 73.800 73.000 74.600 ;
        RECT 74.300 74.400 74.700 74.800 ;
        RECT 75.200 74.900 75.500 75.900 ;
        RECT 75.200 74.500 75.700 74.900 ;
        RECT 75.200 73.700 75.500 74.500 ;
        RECT 76.000 74.200 76.300 75.900 ;
        RECT 77.400 74.800 77.900 75.200 ;
        RECT 77.500 74.400 77.900 74.800 ;
        RECT 78.400 74.900 78.700 75.900 ;
        RECT 78.400 74.500 78.900 74.900 ;
        RECT 75.800 73.800 76.300 74.200 ;
        RECT 69.400 72.800 71.400 73.100 ;
        RECT 69.900 71.100 70.300 72.800 ;
        RECT 71.100 72.400 71.500 72.800 ;
        RECT 71.800 71.100 72.200 73.100 ;
        RECT 74.200 73.400 75.500 73.700 ;
        RECT 74.200 71.100 74.600 73.400 ;
        RECT 76.000 73.100 76.300 73.800 ;
        RECT 78.400 73.700 78.700 74.500 ;
        RECT 79.200 74.200 79.500 75.900 ;
        RECT 80.600 74.800 81.100 75.200 ;
        RECT 80.700 74.400 81.100 74.800 ;
        RECT 81.600 74.900 81.900 75.900 ;
        RECT 81.600 74.500 82.100 74.900 ;
        RECT 79.000 74.100 79.500 74.200 ;
        RECT 79.800 74.100 80.200 74.200 ;
        RECT 79.000 73.800 80.200 74.100 ;
        RECT 75.800 72.800 76.300 73.100 ;
        RECT 77.400 73.400 78.700 73.700 ;
        RECT 75.800 71.100 76.200 72.800 ;
        RECT 77.400 71.100 77.800 73.400 ;
        RECT 79.200 73.100 79.500 73.800 ;
        RECT 81.600 73.700 81.900 74.500 ;
        RECT 82.400 74.200 82.700 75.900 ;
        RECT 82.200 74.100 82.700 74.200 ;
        RECT 83.800 74.100 84.200 74.200 ;
        RECT 82.200 73.800 84.200 74.100 ;
        RECT 79.000 72.800 79.500 73.100 ;
        RECT 80.600 73.400 81.900 73.700 ;
        RECT 79.000 71.100 79.400 72.800 ;
        RECT 80.600 71.100 81.000 73.400 ;
        RECT 82.400 73.100 82.700 73.800 ;
        RECT 83.800 73.400 84.200 73.800 ;
        RECT 82.200 72.800 82.700 73.100 ;
        RECT 84.600 73.100 85.000 79.900 ;
        RECT 85.400 75.800 85.800 76.600 ;
        RECT 86.200 76.200 86.600 79.900 ;
        RECT 87.800 79.600 89.800 79.900 ;
        RECT 87.800 76.200 88.200 79.600 ;
        RECT 86.200 75.900 88.200 76.200 ;
        RECT 88.600 75.900 89.000 79.300 ;
        RECT 89.400 75.900 89.800 79.600 ;
        RECT 88.600 75.600 88.900 75.900 ;
        RECT 86.600 75.200 87.000 75.400 ;
        RECT 87.900 75.300 88.900 75.600 ;
        RECT 87.900 75.200 88.200 75.300 ;
        RECT 86.200 74.900 87.000 75.200 ;
        RECT 86.200 74.800 86.600 74.900 ;
        RECT 87.800 74.800 88.200 75.200 ;
        RECT 89.400 74.800 89.800 75.600 ;
        RECT 85.400 74.100 85.800 74.200 ;
        RECT 87.000 74.100 87.400 74.600 ;
        RECT 85.400 73.800 87.400 74.100 ;
        RECT 87.900 73.100 88.200 74.800 ;
        RECT 88.500 74.400 88.900 74.800 ;
        RECT 88.600 74.200 88.900 74.400 ;
        RECT 88.600 73.800 89.000 74.200 ;
        RECT 90.200 73.400 90.600 74.200 ;
        RECT 91.000 73.200 91.400 79.900 ;
        RECT 92.600 79.600 94.600 79.900 ;
        RECT 91.800 75.800 92.200 76.600 ;
        RECT 92.600 75.900 93.000 79.600 ;
        RECT 93.400 75.900 93.800 79.300 ;
        RECT 94.200 76.200 94.600 79.600 ;
        RECT 95.800 76.200 96.200 79.900 ;
        RECT 94.200 75.900 96.200 76.200 ;
        RECT 96.600 76.200 97.000 79.900 ;
        RECT 98.200 76.200 98.600 79.900 ;
        RECT 96.600 75.900 98.600 76.200 ;
        RECT 99.000 75.900 99.400 79.900 ;
        RECT 101.400 76.200 101.800 79.900 ;
        RECT 103.000 76.200 103.400 79.900 ;
        RECT 101.400 75.900 103.400 76.200 ;
        RECT 103.800 75.900 104.200 79.900 ;
        RECT 93.500 75.600 93.800 75.900 ;
        RECT 92.600 74.800 93.000 75.600 ;
        RECT 93.500 75.300 94.500 75.600 ;
        RECT 94.200 75.200 94.500 75.300 ;
        RECT 95.400 75.200 95.800 75.400 ;
        RECT 97.000 75.200 97.400 75.400 ;
        RECT 99.000 75.200 99.300 75.900 ;
        RECT 101.800 75.200 102.200 75.400 ;
        RECT 103.800 75.200 104.100 75.900 ;
        RECT 94.200 74.800 94.600 75.200 ;
        RECT 95.400 74.900 96.200 75.200 ;
        RECT 95.800 74.800 96.200 74.900 ;
        RECT 96.600 74.900 97.400 75.200 ;
        RECT 98.200 74.900 99.400 75.200 ;
        RECT 96.600 74.800 97.000 74.900 ;
        RECT 93.500 74.400 93.900 74.800 ;
        RECT 93.500 74.200 93.800 74.400 ;
        RECT 91.800 74.100 92.200 74.200 ;
        RECT 93.400 74.100 93.800 74.200 ;
        RECT 91.800 73.800 93.800 74.100 ;
        RECT 84.600 72.800 85.500 73.100 ;
        RECT 82.200 71.100 82.600 72.800 ;
        RECT 85.100 72.200 85.500 72.800 ;
        RECT 85.100 71.800 85.800 72.200 ;
        RECT 85.100 71.100 85.500 71.800 ;
        RECT 87.700 71.100 88.500 73.100 ;
        RECT 91.000 72.800 92.200 73.200 ;
        RECT 94.200 73.100 94.500 74.800 ;
        RECT 95.000 74.100 95.400 74.600 ;
        RECT 97.400 74.100 97.800 74.600 ;
        RECT 95.000 73.800 97.800 74.100 ;
        RECT 98.200 73.100 98.500 74.900 ;
        RECT 99.000 74.800 99.400 74.900 ;
        RECT 101.400 74.900 102.200 75.200 ;
        RECT 103.000 74.900 104.200 75.200 ;
        RECT 101.400 74.800 101.800 74.900 ;
        RECT 102.200 73.800 102.600 74.600 ;
        RECT 91.500 71.100 91.900 72.800 ;
        RECT 93.900 71.100 94.700 73.100 ;
        RECT 98.200 71.100 98.600 73.100 ;
        RECT 99.000 72.800 99.400 73.200 ;
        RECT 103.000 73.100 103.300 74.900 ;
        RECT 103.800 74.800 104.200 74.900 ;
        RECT 103.800 74.100 104.200 74.200 ;
        RECT 104.600 74.100 105.000 74.200 ;
        RECT 103.800 73.800 105.000 74.100 ;
        RECT 104.600 73.400 105.000 73.800 ;
        RECT 98.900 72.400 99.300 72.800 ;
        RECT 103.000 71.100 103.400 73.100 ;
        RECT 103.800 72.800 104.200 73.200 ;
        RECT 105.400 73.100 105.800 79.900 ;
        RECT 106.200 75.800 106.600 77.200 ;
        RECT 108.300 76.300 108.700 79.900 ;
        RECT 107.800 75.900 108.700 76.300 ;
        RECT 107.900 74.200 108.200 75.900 ;
        RECT 108.600 74.800 109.000 75.600 ;
        RECT 107.800 73.800 108.200 74.200 ;
        RECT 105.400 72.800 106.300 73.100 ;
        RECT 103.700 72.400 104.100 72.800 ;
        RECT 105.900 71.100 106.300 72.800 ;
        RECT 107.000 72.400 107.400 73.200 ;
        RECT 107.900 72.200 108.200 73.800 ;
        RECT 109.400 73.400 109.800 74.200 ;
        RECT 110.200 73.100 110.600 79.900 ;
        RECT 111.800 77.900 112.200 79.900 ;
        RECT 111.900 77.800 112.200 77.900 ;
        RECT 113.400 77.900 113.800 79.900 ;
        RECT 115.000 77.900 115.400 79.900 ;
        RECT 113.400 77.800 113.700 77.900 ;
        RECT 111.900 77.500 113.700 77.800 ;
        RECT 115.100 77.800 115.400 77.900 ;
        RECT 116.600 77.900 117.000 79.900 ;
        RECT 116.600 77.800 116.900 77.900 ;
        RECT 115.100 77.500 116.900 77.800 ;
        RECT 111.000 75.800 111.400 76.600 ;
        RECT 111.900 76.200 112.200 77.500 ;
        RECT 112.600 76.400 113.000 77.200 ;
        RECT 115.100 76.200 115.400 77.500 ;
        RECT 115.800 76.400 116.200 77.200 ;
        RECT 111.800 75.800 112.200 76.200 ;
        RECT 111.900 74.200 112.200 75.800 ;
        RECT 114.200 75.400 114.600 76.200 ;
        RECT 115.000 75.800 115.400 76.200 ;
        RECT 113.000 74.800 113.800 75.200 ;
        RECT 115.100 74.200 115.400 75.800 ;
        RECT 117.400 76.100 117.800 76.200 ;
        RECT 118.200 76.100 118.600 79.900 ;
        RECT 120.600 77.900 121.000 79.900 ;
        RECT 120.700 77.800 121.000 77.900 ;
        RECT 122.200 77.900 122.600 79.900 ;
        RECT 122.200 77.800 122.500 77.900 ;
        RECT 120.700 77.500 122.500 77.800 ;
        RECT 121.400 76.400 121.800 77.200 ;
        RECT 122.200 76.200 122.500 77.500 ;
        RECT 123.000 76.200 123.400 79.900 ;
        RECT 124.600 76.200 125.000 79.900 ;
        RECT 117.400 75.800 118.600 76.100 ;
        RECT 117.400 75.400 117.800 75.800 ;
        RECT 116.200 74.800 117.000 75.200 ;
        RECT 111.900 73.900 113.000 74.200 ;
        RECT 115.100 74.100 115.900 74.200 ;
        RECT 115.100 73.900 116.000 74.100 ;
        RECT 112.400 73.800 113.000 73.900 ;
        RECT 110.200 72.800 111.100 73.100 ;
        RECT 107.800 71.100 108.200 72.200 ;
        RECT 110.700 72.200 111.100 72.800 ;
        RECT 110.700 71.800 111.400 72.200 ;
        RECT 110.700 71.100 111.100 71.800 ;
        RECT 112.400 71.100 112.800 73.800 ;
        RECT 115.600 72.200 116.000 73.900 ;
        RECT 115.600 71.800 116.200 72.200 ;
        RECT 115.600 71.100 116.000 71.800 ;
        RECT 118.200 71.100 118.600 75.800 ;
        RECT 119.800 75.400 120.200 76.200 ;
        RECT 122.200 75.800 122.600 76.200 ;
        RECT 123.000 75.900 125.000 76.200 ;
        RECT 125.400 75.900 125.800 79.900 ;
        RECT 127.000 77.900 127.400 79.900 ;
        RECT 127.100 77.800 127.400 77.900 ;
        RECT 128.600 77.900 129.000 79.900 ;
        RECT 130.700 79.200 131.100 79.900 ;
        RECT 130.200 78.800 131.100 79.200 ;
        RECT 128.600 77.800 128.900 77.900 ;
        RECT 127.100 77.500 128.900 77.800 ;
        RECT 127.800 76.400 128.200 77.200 ;
        RECT 128.600 76.200 128.900 77.500 ;
        RECT 130.700 76.200 131.100 78.800 ;
        RECT 131.400 76.800 131.800 77.200 ;
        RECT 131.500 76.200 131.800 76.800 ;
        RECT 132.600 76.200 133.000 79.900 ;
        RECT 133.300 76.200 133.700 76.300 ;
        RECT 120.600 74.800 121.400 75.200 ;
        RECT 122.200 74.200 122.500 75.800 ;
        RECT 123.400 75.200 123.800 75.400 ;
        RECT 125.400 75.200 125.700 75.900 ;
        RECT 126.200 75.400 126.600 76.200 ;
        RECT 128.600 75.800 129.000 76.200 ;
        RECT 130.700 75.900 131.200 76.200 ;
        RECT 131.500 75.900 132.200 76.200 ;
        RECT 132.600 75.900 133.700 76.200 ;
        RECT 134.800 76.200 135.600 79.900 ;
        RECT 136.600 76.200 137.000 76.300 ;
        RECT 137.400 76.200 137.800 79.900 ;
        RECT 139.000 77.800 139.400 79.900 ;
        RECT 140.600 77.900 141.000 79.900 ;
        RECT 142.200 77.900 142.600 79.900 ;
        RECT 140.600 77.800 140.900 77.900 ;
        RECT 139.100 77.500 140.900 77.800 ;
        RECT 142.300 77.800 142.600 77.900 ;
        RECT 143.800 77.900 144.200 79.900 ;
        RECT 144.600 77.900 145.000 79.900 ;
        RECT 143.800 77.800 144.100 77.900 ;
        RECT 142.300 77.500 144.100 77.800 ;
        RECT 134.800 75.900 135.800 76.200 ;
        RECT 136.600 75.900 137.800 76.200 ;
        RECT 138.200 76.800 138.600 77.200 ;
        RECT 138.200 76.200 138.500 76.800 ;
        RECT 139.800 76.400 140.200 77.200 ;
        RECT 140.600 76.200 140.900 77.500 ;
        RECT 141.400 77.100 141.800 77.200 ;
        RECT 143.000 77.100 143.400 77.200 ;
        RECT 141.400 76.800 143.400 77.100 ;
        RECT 143.000 76.400 143.400 76.800 ;
        RECT 143.800 76.200 144.100 77.500 ;
        RECT 144.700 77.800 145.000 77.900 ;
        RECT 146.200 77.900 146.600 79.900 ;
        RECT 146.200 77.800 146.500 77.900 ;
        RECT 144.700 77.500 146.500 77.800 ;
        RECT 144.700 76.200 145.000 77.500 ;
        RECT 145.400 76.400 145.800 77.200 ;
        RECT 147.800 76.200 148.200 79.900 ;
        RECT 149.400 76.200 149.800 79.900 ;
        RECT 123.000 74.900 123.800 75.200 ;
        RECT 124.600 74.900 125.800 75.200 ;
        RECT 123.000 74.800 123.400 74.900 ;
        RECT 119.000 73.400 119.400 74.200 ;
        RECT 121.700 74.100 122.500 74.200 ;
        RECT 121.600 73.900 122.500 74.100 ;
        RECT 121.600 72.200 122.000 73.900 ;
        RECT 123.800 73.800 124.200 74.600 ;
        RECT 124.600 74.100 124.900 74.900 ;
        RECT 125.400 74.800 125.800 74.900 ;
        RECT 127.000 74.800 127.800 75.200 ;
        RECT 128.600 74.200 128.900 75.800 ;
        RECT 130.200 74.400 130.600 75.200 ;
        RECT 130.900 74.200 131.200 75.900 ;
        RECT 131.800 75.800 132.200 75.900 ;
        RECT 133.400 75.600 133.700 75.900 ;
        RECT 133.400 75.300 135.100 75.600 ;
        RECT 134.700 75.200 135.100 75.300 ;
        RECT 135.500 75.200 135.800 75.900 ;
        RECT 135.500 75.100 136.200 75.200 ;
        RECT 138.200 75.100 138.600 76.200 ;
        RECT 140.600 75.800 141.000 76.200 ;
        RECT 133.600 74.900 134.000 75.000 ;
        RECT 135.500 74.900 138.600 75.100 ;
        RECT 133.600 74.600 134.900 74.900 ;
        RECT 134.600 74.300 134.900 74.600 ;
        RECT 135.300 74.800 138.600 74.900 ;
        RECT 139.000 74.800 139.800 75.200 ;
        RECT 135.300 74.600 135.800 74.800 ;
        RECT 125.400 74.100 125.800 74.200 ;
        RECT 128.100 74.100 128.900 74.200 ;
        RECT 124.600 73.800 125.800 74.100 ;
        RECT 128.000 73.900 128.900 74.100 ;
        RECT 129.400 74.100 129.800 74.200 ;
        RECT 121.400 71.800 122.000 72.200 ;
        RECT 121.600 71.100 122.000 71.800 ;
        RECT 124.600 73.100 124.900 73.800 ;
        RECT 124.600 71.100 125.000 73.100 ;
        RECT 125.400 72.800 125.800 73.200 ;
        RECT 125.300 72.400 125.700 72.800 ;
        RECT 128.000 71.100 128.400 73.900 ;
        RECT 129.400 73.800 130.200 74.100 ;
        RECT 130.900 73.800 132.200 74.200 ;
        RECT 132.600 74.100 133.400 74.200 ;
        RECT 132.600 73.800 134.300 74.100 ;
        RECT 134.600 73.900 135.000 74.300 ;
        RECT 129.800 73.600 130.200 73.800 ;
        RECT 129.500 73.100 131.300 73.300 ;
        RECT 131.800 73.100 132.100 73.800 ;
        RECT 134.000 73.600 134.300 73.800 ;
        RECT 133.300 73.400 133.700 73.500 ;
        RECT 132.600 73.100 133.700 73.400 ;
        RECT 134.000 73.300 135.000 73.600 ;
        RECT 134.200 73.200 135.000 73.300 ;
        RECT 129.400 73.000 131.400 73.100 ;
        RECT 129.400 71.100 129.800 73.000 ;
        RECT 131.000 71.100 131.400 73.000 ;
        RECT 131.800 71.100 132.200 73.100 ;
        RECT 132.600 71.100 133.000 73.100 ;
        RECT 135.300 72.900 135.600 74.600 ;
        RECT 140.600 74.200 140.900 75.800 ;
        RECT 141.400 75.400 141.800 76.200 ;
        RECT 143.800 75.800 144.200 76.200 ;
        RECT 144.600 75.800 145.000 76.200 ;
        RECT 142.200 74.800 143.000 75.200 ;
        RECT 143.800 74.200 144.100 75.800 ;
        RECT 136.000 73.800 136.400 74.200 ;
        RECT 137.000 73.800 137.800 74.200 ;
        RECT 140.100 74.100 140.900 74.200 ;
        RECT 143.300 74.100 144.100 74.200 ;
        RECT 140.000 73.900 140.900 74.100 ;
        RECT 143.200 73.900 144.100 74.100 ;
        RECT 144.700 74.200 145.000 75.800 ;
        RECT 147.000 75.400 147.400 76.200 ;
        RECT 147.800 75.900 149.800 76.200 ;
        RECT 150.200 75.900 150.600 79.900 ;
        RECT 148.200 75.200 148.600 75.400 ;
        RECT 150.200 75.200 150.500 75.900 ;
        RECT 145.800 74.800 146.600 75.200 ;
        RECT 147.800 74.900 148.600 75.200 ;
        RECT 149.400 74.900 150.600 75.200 ;
        RECT 147.800 74.800 148.200 74.900 ;
        RECT 144.700 74.100 145.500 74.200 ;
        RECT 144.700 73.900 145.600 74.100 ;
        RECT 136.000 73.600 136.300 73.800 ;
        RECT 135.900 73.200 136.300 73.600 ;
        RECT 136.600 73.400 137.000 73.500 ;
        RECT 136.600 73.100 137.800 73.400 ;
        RECT 134.800 71.100 135.600 72.900 ;
        RECT 137.400 71.100 137.800 73.100 ;
        RECT 140.000 71.100 140.400 73.900 ;
        RECT 143.200 72.200 143.600 73.900 ;
        RECT 145.200 72.200 145.600 73.900 ;
        RECT 148.600 73.800 149.000 74.600 ;
        RECT 149.400 73.100 149.700 74.900 ;
        RECT 150.200 74.800 150.600 74.900 ;
        RECT 143.200 71.800 144.200 72.200 ;
        RECT 145.200 71.800 145.800 72.200 ;
        RECT 143.200 71.100 143.600 71.800 ;
        RECT 145.200 71.100 145.600 71.800 ;
        RECT 149.400 71.100 149.800 73.100 ;
        RECT 150.200 72.800 150.600 73.200 ;
        RECT 150.100 72.400 150.500 72.800 ;
        RECT 1.400 68.900 1.800 69.900 ;
        RECT 1.500 67.200 1.800 68.900 ;
        RECT 1.400 67.100 1.800 67.200 ;
        RECT 2.200 67.800 2.600 68.200 ;
        RECT 3.000 67.900 3.400 69.900 ;
        RECT 5.200 68.100 6.000 69.900 ;
        RECT 2.200 67.100 2.500 67.800 ;
        RECT 3.000 67.600 4.200 67.900 ;
        RECT 3.800 67.500 4.200 67.600 ;
        RECT 1.400 66.800 2.500 67.100 ;
        RECT 1.500 65.100 1.800 66.800 ;
        RECT 5.200 66.400 5.500 68.100 ;
        RECT 7.800 67.900 8.200 69.900 ;
        RECT 7.100 67.600 8.200 67.900 ;
        RECT 8.600 67.800 9.000 68.600 ;
        RECT 7.100 67.500 7.500 67.600 ;
        RECT 5.800 66.700 6.200 67.100 ;
        RECT 5.000 66.200 5.500 66.400 ;
        RECT 4.600 66.100 5.500 66.200 ;
        RECT 5.900 66.400 6.200 66.700 ;
        RECT 5.900 66.100 7.200 66.400 ;
        RECT 4.600 65.800 5.300 66.100 ;
        RECT 6.800 66.000 7.200 66.100 ;
        RECT 9.400 66.100 9.800 69.900 ;
        RECT 11.800 67.900 12.200 69.900 ;
        RECT 14.200 68.900 14.600 69.900 ;
        RECT 16.100 69.200 16.500 69.900 ;
        RECT 12.500 68.200 12.900 68.600 ;
        RECT 11.000 66.400 11.400 67.200 ;
        RECT 10.200 66.100 10.600 66.200 ;
        RECT 11.800 66.100 12.100 67.900 ;
        RECT 12.600 67.800 13.000 68.200 ;
        RECT 14.200 67.200 14.500 68.900 ;
        RECT 15.800 68.800 16.500 69.200 ;
        RECT 15.000 67.800 15.400 68.600 ;
        RECT 16.100 68.200 16.500 68.800 ;
        RECT 16.100 67.900 17.000 68.200 ;
        RECT 14.200 66.800 14.600 67.200 ;
        RECT 15.800 66.800 16.200 67.200 ;
        RECT 12.600 66.100 13.000 66.200 ;
        RECT 9.400 65.800 11.000 66.100 ;
        RECT 11.800 65.800 13.000 66.100 ;
        RECT 5.000 65.100 5.300 65.800 ;
        RECT 5.700 65.700 6.100 65.800 ;
        RECT 5.700 65.400 7.400 65.700 ;
        RECT 7.100 65.100 7.400 65.400 ;
        RECT 1.400 64.700 2.300 65.100 ;
        RECT 1.900 61.100 2.300 64.700 ;
        RECT 3.000 64.800 4.200 65.100 ;
        RECT 5.000 64.800 6.000 65.100 ;
        RECT 3.000 61.100 3.400 64.800 ;
        RECT 3.800 64.700 4.200 64.800 ;
        RECT 5.200 61.100 6.000 64.800 ;
        RECT 7.100 64.800 8.200 65.100 ;
        RECT 7.100 64.700 7.500 64.800 ;
        RECT 7.800 61.100 8.200 64.800 ;
        RECT 9.400 61.100 9.800 65.800 ;
        RECT 10.600 65.600 11.000 65.800 ;
        RECT 12.600 65.100 12.900 65.800 ;
        RECT 13.400 65.400 13.800 66.200 ;
        RECT 14.200 66.100 14.500 66.800 ;
        RECT 15.800 66.100 16.100 66.800 ;
        RECT 14.200 65.800 16.100 66.100 ;
        RECT 14.200 65.100 14.500 65.800 ;
        RECT 10.200 64.800 12.200 65.100 ;
        RECT 10.200 61.100 10.600 64.800 ;
        RECT 11.800 61.100 12.200 64.800 ;
        RECT 12.600 61.100 13.000 65.100 ;
        RECT 13.700 64.700 14.600 65.100 ;
        RECT 13.700 61.100 14.100 64.700 ;
        RECT 15.800 64.400 16.200 65.200 ;
        RECT 16.600 61.100 17.000 67.900 ;
        RECT 18.200 67.900 18.600 69.900 ;
        RECT 20.400 69.200 21.200 69.900 ;
        RECT 20.400 68.800 21.800 69.200 ;
        RECT 20.400 68.100 21.200 68.800 ;
        RECT 18.200 67.600 19.400 67.900 ;
        RECT 17.400 67.100 17.800 67.600 ;
        RECT 19.000 67.500 19.400 67.600 ;
        RECT 19.700 67.400 20.100 67.800 ;
        RECT 19.700 67.200 20.000 67.400 ;
        RECT 18.200 67.100 19.000 67.200 ;
        RECT 17.400 66.800 19.000 67.100 ;
        RECT 19.600 66.800 20.000 67.200 ;
        RECT 20.400 67.100 20.700 68.100 ;
        RECT 23.000 67.900 23.400 69.900 ;
        RECT 21.000 67.400 21.800 67.800 ;
        RECT 22.100 67.600 23.400 67.900 ;
        RECT 23.800 67.900 24.200 69.900 ;
        RECT 26.000 69.200 26.800 69.900 ;
        RECT 26.000 68.800 27.400 69.200 ;
        RECT 26.000 68.100 26.800 68.800 ;
        RECT 23.800 67.600 25.000 67.900 ;
        RECT 22.100 67.500 22.500 67.600 ;
        RECT 24.600 67.500 25.000 67.600 ;
        RECT 25.300 67.400 25.700 67.800 ;
        RECT 25.300 67.200 25.600 67.400 ;
        RECT 22.600 67.100 23.400 67.200 ;
        RECT 20.400 66.800 20.900 67.100 ;
        RECT 22.300 67.000 23.400 67.100 ;
        RECT 20.600 66.200 20.900 66.800 ;
        RECT 21.200 66.800 23.400 67.000 ;
        RECT 23.800 66.800 24.600 67.200 ;
        RECT 25.200 66.800 25.600 67.200 ;
        RECT 26.000 67.100 26.300 68.100 ;
        RECT 28.600 67.900 29.000 69.900 ;
        RECT 26.600 67.400 27.400 67.800 ;
        RECT 27.700 67.600 29.000 67.900 ;
        RECT 29.400 67.900 29.800 69.900 ;
        RECT 31.600 68.100 32.400 69.900 ;
        RECT 29.400 67.600 30.600 67.900 ;
        RECT 27.700 67.500 28.100 67.600 ;
        RECT 30.200 67.500 30.600 67.600 ;
        RECT 30.900 67.400 31.300 67.800 ;
        RECT 30.900 67.200 31.200 67.400 ;
        RECT 28.200 67.100 29.000 67.200 ;
        RECT 26.000 66.800 26.500 67.100 ;
        RECT 27.900 67.000 29.000 67.100 ;
        RECT 21.200 66.700 22.600 66.800 ;
        RECT 21.200 66.600 21.600 66.700 ;
        RECT 26.200 66.200 26.500 66.800 ;
        RECT 26.800 66.800 29.000 67.000 ;
        RECT 29.400 66.800 30.200 67.200 ;
        RECT 30.800 66.800 31.200 67.200 ;
        RECT 31.600 67.100 31.900 68.100 ;
        RECT 34.200 67.900 34.600 69.900 ;
        RECT 35.800 68.900 36.200 69.900 ;
        RECT 32.200 67.400 33.000 67.800 ;
        RECT 33.300 67.600 34.600 67.900 ;
        RECT 35.000 67.800 35.400 68.600 ;
        RECT 33.300 67.500 33.700 67.600 ;
        RECT 35.900 67.200 36.200 68.900 ;
        RECT 37.400 67.500 37.800 69.900 ;
        RECT 39.600 69.200 40.000 69.900 ;
        RECT 39.000 68.900 40.000 69.200 ;
        RECT 41.800 68.900 42.200 69.900 ;
        RECT 43.900 69.200 44.500 69.900 ;
        RECT 43.800 68.900 44.500 69.200 ;
        RECT 39.000 68.500 39.400 68.900 ;
        RECT 41.800 68.600 42.100 68.900 ;
        RECT 39.800 68.200 40.200 68.600 ;
        RECT 40.700 68.300 42.100 68.600 ;
        RECT 43.800 68.500 44.200 68.900 ;
        RECT 40.700 68.200 41.100 68.300 ;
        RECT 33.800 67.100 34.600 67.200 ;
        RECT 35.800 67.100 36.200 67.200 ;
        RECT 31.600 66.800 32.100 67.100 ;
        RECT 33.500 67.000 36.200 67.100 ;
        RECT 26.800 66.700 28.200 66.800 ;
        RECT 26.800 66.600 27.200 66.700 ;
        RECT 31.800 66.200 32.100 66.800 ;
        RECT 32.400 66.800 36.200 67.000 ;
        RECT 37.800 67.100 38.600 67.200 ;
        RECT 39.900 67.100 40.200 68.200 ;
        RECT 44.700 67.700 45.100 67.800 ;
        RECT 46.200 67.700 46.600 69.900 ;
        RECT 44.700 67.400 46.600 67.700 ;
        RECT 48.600 67.500 49.000 69.900 ;
        RECT 50.800 69.200 51.200 69.900 ;
        RECT 50.200 68.900 51.200 69.200 ;
        RECT 53.000 68.900 53.400 69.900 ;
        RECT 55.100 69.200 55.700 69.900 ;
        RECT 55.000 68.900 55.700 69.200 ;
        RECT 50.200 68.500 50.600 68.900 ;
        RECT 53.000 68.600 53.300 68.900 ;
        RECT 51.000 68.200 51.400 68.600 ;
        RECT 51.900 68.300 53.300 68.600 ;
        RECT 55.000 68.500 55.400 68.900 ;
        RECT 51.900 68.200 52.300 68.300 ;
        RECT 42.700 67.100 43.100 67.200 ;
        RECT 37.800 66.800 43.300 67.100 ;
        RECT 32.400 66.700 33.800 66.800 ;
        RECT 32.400 66.600 32.800 66.700 ;
        RECT 20.600 65.800 21.000 66.200 ;
        RECT 21.900 66.100 22.300 66.200 ;
        RECT 21.500 65.800 22.300 66.100 ;
        RECT 26.200 65.800 26.600 66.200 ;
        RECT 27.500 66.100 27.900 66.200 ;
        RECT 27.100 65.800 27.900 66.100 ;
        RECT 31.000 66.100 31.400 66.200 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 33.100 66.100 33.500 66.200 ;
        RECT 31.000 65.800 32.200 66.100 ;
        RECT 32.700 65.800 33.500 66.100 ;
        RECT 20.600 65.100 20.900 65.800 ;
        RECT 21.500 65.700 21.900 65.800 ;
        RECT 26.200 65.100 26.500 65.800 ;
        RECT 27.100 65.700 27.500 65.800 ;
        RECT 31.800 65.100 32.100 65.800 ;
        RECT 32.700 65.700 33.100 65.800 ;
        RECT 35.900 65.100 36.200 66.800 ;
        RECT 39.300 66.700 39.700 66.800 ;
        RECT 38.500 66.200 38.900 66.300 ;
        RECT 39.800 66.200 40.200 66.300 ;
        RECT 43.000 66.200 43.300 66.800 ;
        RECT 43.800 66.400 44.200 66.500 ;
        RECT 36.600 65.400 37.000 66.200 ;
        RECT 38.500 65.900 41.000 66.200 ;
        RECT 40.600 65.800 41.000 65.900 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 43.800 66.100 45.700 66.400 ;
        RECT 45.300 66.000 45.700 66.100 ;
        RECT 37.400 65.500 40.200 65.600 ;
        RECT 37.400 65.400 40.300 65.500 ;
        RECT 37.400 65.300 42.300 65.400 ;
        RECT 18.200 64.800 19.400 65.100 ;
        RECT 18.200 61.100 18.600 64.800 ;
        RECT 19.000 64.700 19.400 64.800 ;
        RECT 20.400 61.100 21.200 65.100 ;
        RECT 22.100 64.800 23.400 65.100 ;
        RECT 22.100 64.700 22.500 64.800 ;
        RECT 23.000 61.100 23.400 64.800 ;
        RECT 23.800 64.800 25.000 65.100 ;
        RECT 23.800 61.100 24.200 64.800 ;
        RECT 24.600 64.700 25.000 64.800 ;
        RECT 26.000 61.100 26.800 65.100 ;
        RECT 27.700 64.800 29.000 65.100 ;
        RECT 27.700 64.700 28.100 64.800 ;
        RECT 28.600 61.100 29.000 64.800 ;
        RECT 29.400 64.800 30.600 65.100 ;
        RECT 29.400 61.100 29.800 64.800 ;
        RECT 30.200 64.700 30.600 64.800 ;
        RECT 31.600 61.100 32.400 65.100 ;
        RECT 33.300 64.800 34.600 65.100 ;
        RECT 33.300 64.700 33.700 64.800 ;
        RECT 34.200 61.100 34.600 64.800 ;
        RECT 35.800 64.700 36.700 65.100 ;
        RECT 36.300 61.100 36.700 64.700 ;
        RECT 37.400 61.100 37.800 65.300 ;
        RECT 39.900 65.100 42.300 65.300 ;
        RECT 39.000 64.500 41.700 64.800 ;
        RECT 39.000 64.400 39.400 64.500 ;
        RECT 41.300 64.400 41.700 64.500 ;
        RECT 42.000 64.500 42.300 65.100 ;
        RECT 43.000 65.200 43.300 65.800 ;
        RECT 44.500 65.700 44.900 65.800 ;
        RECT 46.200 65.700 46.600 67.400 ;
        RECT 49.000 67.100 49.800 67.200 ;
        RECT 51.100 67.100 51.400 68.200 ;
        RECT 55.900 67.700 56.300 67.800 ;
        RECT 57.400 67.700 57.800 69.900 ;
        RECT 59.500 69.200 59.900 69.900 ;
        RECT 59.500 68.800 60.200 69.200 ;
        RECT 59.500 68.200 59.900 68.800 ;
        RECT 61.900 68.200 62.300 69.900 ;
        RECT 55.900 67.400 57.800 67.700 ;
        RECT 59.000 67.900 59.900 68.200 ;
        RECT 61.400 67.900 62.300 68.200 ;
        RECT 52.600 67.100 53.000 67.200 ;
        RECT 53.900 67.100 54.300 67.200 ;
        RECT 49.000 66.800 54.500 67.100 ;
        RECT 50.500 66.700 50.900 66.800 ;
        RECT 49.700 66.200 50.100 66.300 ;
        RECT 51.000 66.200 51.400 66.300 ;
        RECT 49.700 65.900 52.200 66.200 ;
        RECT 51.800 65.800 52.200 65.900 ;
        RECT 44.500 65.400 46.600 65.700 ;
        RECT 43.000 64.900 44.200 65.200 ;
        RECT 42.700 64.500 43.100 64.600 ;
        RECT 42.000 64.200 43.100 64.500 ;
        RECT 43.900 64.400 44.200 64.900 ;
        RECT 43.900 64.000 44.600 64.400 ;
        RECT 40.700 63.700 41.100 63.800 ;
        RECT 42.100 63.700 42.500 63.800 ;
        RECT 39.000 63.100 39.400 63.500 ;
        RECT 40.700 63.400 42.500 63.700 ;
        RECT 41.800 63.100 42.100 63.400 ;
        RECT 43.800 63.100 44.200 63.500 ;
        RECT 39.000 62.800 40.000 63.100 ;
        RECT 39.600 61.100 40.000 62.800 ;
        RECT 41.800 61.100 42.200 63.100 ;
        RECT 43.900 61.100 44.500 63.100 ;
        RECT 46.200 61.100 46.600 65.400 ;
        RECT 48.600 65.500 51.400 65.600 ;
        RECT 48.600 65.400 51.500 65.500 ;
        RECT 48.600 65.300 53.500 65.400 ;
        RECT 48.600 61.100 49.000 65.300 ;
        RECT 51.100 65.100 53.500 65.300 ;
        RECT 50.200 64.500 52.900 64.800 ;
        RECT 50.200 64.400 50.600 64.500 ;
        RECT 52.500 64.400 52.900 64.500 ;
        RECT 53.200 64.500 53.500 65.100 ;
        RECT 54.200 65.200 54.500 66.800 ;
        RECT 55.000 66.400 55.400 66.500 ;
        RECT 55.000 66.100 56.900 66.400 ;
        RECT 56.500 66.000 56.900 66.100 ;
        RECT 55.700 65.700 56.100 65.800 ;
        RECT 57.400 65.700 57.800 67.400 ;
        RECT 58.200 66.800 58.600 67.600 ;
        RECT 55.700 65.400 57.800 65.700 ;
        RECT 54.200 64.900 55.400 65.200 ;
        RECT 53.900 64.500 54.300 64.600 ;
        RECT 53.200 64.200 54.300 64.500 ;
        RECT 55.100 64.400 55.400 64.900 ;
        RECT 55.100 64.000 55.800 64.400 ;
        RECT 51.900 63.700 52.300 63.800 ;
        RECT 53.300 63.700 53.700 63.800 ;
        RECT 50.200 63.100 50.600 63.500 ;
        RECT 51.900 63.400 53.700 63.700 ;
        RECT 53.000 63.100 53.300 63.400 ;
        RECT 55.000 63.100 55.400 63.500 ;
        RECT 50.200 62.800 51.200 63.100 ;
        RECT 50.800 61.100 51.200 62.800 ;
        RECT 53.000 61.100 53.400 63.100 ;
        RECT 55.100 61.100 55.700 63.100 ;
        RECT 57.400 61.100 57.800 65.400 ;
        RECT 59.000 61.100 59.400 67.900 ;
        RECT 60.600 66.800 61.000 67.600 ;
        RECT 61.400 66.100 61.800 67.900 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 63.600 67.100 64.000 69.900 ;
        RECT 66.800 68.100 67.200 69.900 ;
        RECT 67.800 68.100 68.200 68.200 ;
        RECT 66.800 67.800 68.200 68.100 ;
        RECT 69.400 67.800 69.800 68.600 ;
        RECT 66.800 67.100 67.200 67.800 ;
        RECT 63.100 66.900 64.000 67.100 ;
        RECT 66.300 66.900 67.200 67.100 ;
        RECT 63.100 66.800 63.900 66.900 ;
        RECT 66.300 66.800 67.100 66.900 ;
        RECT 62.200 66.100 62.500 66.800 ;
        RECT 61.400 65.800 62.500 66.100 ;
        RECT 59.800 65.100 60.200 65.200 ;
        RECT 60.600 65.100 61.000 65.200 ;
        RECT 59.800 64.800 61.000 65.100 ;
        RECT 59.800 64.400 60.200 64.800 ;
        RECT 61.400 61.100 61.800 65.800 ;
        RECT 63.100 65.200 63.400 66.800 ;
        RECT 64.200 65.800 65.000 66.200 ;
        RECT 62.200 64.400 62.600 65.200 ;
        RECT 63.000 64.800 63.400 65.200 ;
        RECT 65.400 64.800 65.800 65.600 ;
        RECT 66.300 65.200 66.600 66.800 ;
        RECT 67.400 65.800 68.200 66.200 ;
        RECT 66.200 64.800 66.600 65.200 ;
        RECT 68.600 65.100 69.000 65.600 ;
        RECT 70.200 65.100 70.600 69.900 ;
        RECT 71.000 67.900 71.400 69.900 ;
        RECT 71.800 68.000 72.200 69.900 ;
        RECT 73.400 68.000 73.800 69.900 ;
        RECT 71.800 67.900 73.800 68.000 ;
        RECT 74.200 68.000 74.600 69.900 ;
        RECT 75.800 68.000 76.200 69.900 ;
        RECT 74.200 67.900 76.200 68.000 ;
        RECT 76.600 67.900 77.000 69.900 ;
        RECT 78.700 68.200 79.100 69.900 ;
        RECT 81.100 68.200 81.500 69.900 ;
        RECT 83.000 68.200 83.400 69.900 ;
        RECT 78.200 67.900 79.100 68.200 ;
        RECT 80.600 67.900 81.500 68.200 ;
        RECT 82.900 67.900 83.400 68.200 ;
        RECT 71.100 67.200 71.400 67.900 ;
        RECT 71.900 67.700 73.700 67.900 ;
        RECT 74.300 67.700 76.100 67.900 ;
        RECT 73.000 67.200 73.400 67.400 ;
        RECT 74.600 67.200 75.000 67.400 ;
        RECT 76.600 67.200 76.900 67.900 ;
        RECT 71.000 66.800 72.300 67.200 ;
        RECT 73.000 67.100 73.800 67.200 ;
        RECT 74.200 67.100 75.000 67.200 ;
        RECT 73.000 66.900 75.000 67.100 ;
        RECT 73.400 66.800 74.600 66.900 ;
        RECT 75.700 66.800 77.000 67.200 ;
        RECT 77.400 66.800 77.800 67.600 ;
        RECT 72.000 66.200 72.300 66.800 ;
        RECT 71.800 65.800 72.300 66.200 ;
        RECT 72.600 66.100 73.000 66.600 ;
        RECT 75.000 66.100 75.400 66.600 ;
        RECT 72.600 65.800 75.400 66.100 ;
        RECT 75.700 66.100 76.000 66.800 ;
        RECT 77.400 66.100 77.800 66.200 ;
        RECT 75.700 65.800 77.800 66.100 ;
        RECT 78.200 66.100 78.600 67.900 ;
        RECT 79.800 66.800 80.200 67.600 ;
        RECT 79.000 66.100 79.400 66.200 ;
        RECT 78.200 65.800 79.400 66.100 ;
        RECT 71.000 65.100 71.400 65.200 ;
        RECT 72.000 65.100 72.300 65.800 ;
        RECT 75.700 65.100 76.000 65.800 ;
        RECT 76.600 65.100 77.000 65.200 ;
        RECT 68.600 64.800 71.700 65.100 ;
        RECT 72.000 64.800 72.500 65.100 ;
        RECT 63.100 63.500 63.400 64.800 ;
        RECT 63.800 63.800 64.200 64.600 ;
        RECT 66.300 63.500 66.600 64.800 ;
        RECT 67.000 63.800 67.400 64.600 ;
        RECT 63.100 63.200 64.900 63.500 ;
        RECT 66.300 63.200 68.100 63.500 ;
        RECT 63.100 63.100 63.400 63.200 ;
        RECT 63.000 61.100 63.400 63.100 ;
        RECT 64.600 61.100 65.000 63.200 ;
        RECT 66.300 63.100 66.600 63.200 ;
        RECT 66.200 61.100 66.600 63.100 ;
        RECT 67.800 63.100 68.100 63.200 ;
        RECT 67.800 61.100 68.200 63.100 ;
        RECT 70.200 61.100 70.600 64.800 ;
        RECT 71.400 64.200 71.700 64.800 ;
        RECT 71.400 63.800 71.800 64.200 ;
        RECT 72.100 61.100 72.500 64.800 ;
        RECT 75.500 64.800 76.000 65.100 ;
        RECT 76.300 64.800 77.000 65.100 ;
        RECT 75.500 61.100 75.900 64.800 ;
        RECT 76.300 64.200 76.600 64.800 ;
        RECT 76.200 63.800 76.600 64.200 ;
        RECT 78.200 61.100 78.600 65.800 ;
        RECT 79.000 64.400 79.400 65.200 ;
        RECT 79.800 64.100 80.200 64.200 ;
        RECT 80.600 64.100 81.000 67.900 ;
        RECT 82.900 67.200 83.200 67.900 ;
        RECT 84.600 67.600 85.000 69.900 ;
        RECT 83.700 67.300 85.000 67.600 ;
        RECT 85.400 67.600 85.800 69.900 ;
        RECT 87.000 68.200 87.400 69.900 ;
        RECT 88.900 68.200 89.300 69.900 ;
        RECT 87.000 67.900 87.500 68.200 ;
        RECT 88.900 67.900 89.800 68.200 ;
        RECT 91.000 68.000 91.400 69.900 ;
        RECT 92.600 69.600 94.600 69.900 ;
        RECT 92.600 68.000 93.000 69.600 ;
        RECT 91.000 67.900 93.000 68.000 ;
        RECT 85.400 67.300 86.700 67.600 ;
        RECT 82.200 67.100 82.600 67.200 ;
        RECT 82.900 67.100 83.400 67.200 ;
        RECT 82.200 66.800 83.400 67.100 ;
        RECT 81.400 64.400 81.800 65.200 ;
        RECT 82.900 65.100 83.200 66.800 ;
        RECT 83.700 66.500 84.000 67.300 ;
        RECT 83.500 66.100 84.000 66.500 ;
        RECT 83.700 65.100 84.000 66.100 ;
        RECT 84.500 66.200 84.900 66.600 ;
        RECT 85.500 66.200 85.900 66.600 ;
        RECT 84.500 66.100 85.000 66.200 ;
        RECT 85.400 66.100 85.900 66.200 ;
        RECT 84.500 65.800 85.900 66.100 ;
        RECT 86.400 66.500 86.700 67.300 ;
        RECT 87.200 67.200 87.500 67.900 ;
        RECT 87.000 66.800 87.500 67.200 ;
        RECT 86.400 66.100 86.900 66.500 ;
        RECT 86.400 65.100 86.700 66.100 ;
        RECT 87.200 65.100 87.500 66.800 ;
        RECT 82.900 64.600 83.400 65.100 ;
        RECT 83.700 64.800 85.000 65.100 ;
        RECT 79.800 63.800 81.000 64.100 ;
        RECT 80.600 61.100 81.000 63.800 ;
        RECT 83.000 61.100 83.400 64.600 ;
        RECT 84.600 61.100 85.000 64.800 ;
        RECT 85.400 64.800 86.700 65.100 ;
        RECT 85.400 61.100 85.800 64.800 ;
        RECT 87.000 64.600 87.500 65.100 ;
        RECT 87.000 61.100 87.400 64.600 ;
        RECT 88.600 64.400 89.000 65.200 ;
        RECT 89.400 65.100 89.800 67.900 ;
        RECT 91.100 67.700 92.900 67.900 ;
        RECT 93.400 67.800 93.800 69.300 ;
        RECT 94.200 67.900 94.600 69.600 ;
        RECT 95.000 67.900 95.400 69.900 ;
        RECT 95.800 68.000 96.200 69.900 ;
        RECT 97.400 68.000 97.800 69.900 ;
        RECT 95.800 67.900 97.800 68.000 ;
        RECT 98.200 68.000 98.600 69.900 ;
        RECT 99.800 68.000 100.200 69.900 ;
        RECT 98.200 67.900 100.200 68.000 ;
        RECT 100.600 67.900 101.000 69.900 ;
        RECT 90.200 66.800 90.600 67.600 ;
        RECT 91.400 67.200 91.800 67.400 ;
        RECT 93.500 67.200 93.800 67.800 ;
        RECT 95.100 67.200 95.400 67.900 ;
        RECT 95.900 67.700 97.700 67.900 ;
        RECT 98.300 67.700 100.100 67.900 ;
        RECT 97.000 67.200 97.400 67.400 ;
        RECT 98.600 67.200 99.000 67.400 ;
        RECT 100.600 67.200 100.900 67.900 ;
        RECT 91.000 66.900 91.800 67.200 ;
        RECT 92.600 66.900 93.800 67.200 ;
        RECT 91.000 66.800 91.400 66.900 ;
        RECT 92.600 66.800 93.000 66.900 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 91.800 65.800 92.200 66.600 ;
        RECT 90.200 65.100 90.500 65.800 ;
        RECT 92.600 65.100 92.900 66.800 ;
        RECT 93.400 65.800 93.800 66.600 ;
        RECT 94.200 66.400 94.600 67.200 ;
        RECT 95.000 66.800 96.300 67.200 ;
        RECT 97.000 67.100 97.800 67.200 ;
        RECT 98.200 67.100 99.000 67.200 ;
        RECT 97.000 66.900 99.000 67.100 ;
        RECT 97.400 66.800 98.600 66.900 ;
        RECT 99.700 66.800 101.000 67.200 ;
        RECT 103.000 66.800 103.400 67.600 ;
        RECT 96.000 66.200 96.300 66.800 ;
        RECT 95.800 65.800 96.300 66.200 ;
        RECT 96.600 66.100 97.000 66.600 ;
        RECT 97.400 66.100 97.800 66.200 ;
        RECT 99.000 66.100 99.400 66.600 ;
        RECT 96.600 65.800 99.400 66.100 ;
        RECT 95.000 65.100 95.400 65.200 ;
        RECT 96.000 65.100 96.300 65.800 ;
        RECT 99.700 65.100 100.000 66.800 ;
        RECT 103.800 66.100 104.200 69.900 ;
        RECT 104.600 67.900 105.000 69.900 ;
        RECT 105.400 68.000 105.800 69.900 ;
        RECT 107.000 68.000 107.400 69.900 ;
        RECT 105.400 67.900 107.400 68.000 ;
        RECT 107.800 68.000 108.200 69.900 ;
        RECT 109.400 68.000 109.800 69.900 ;
        RECT 107.800 67.900 109.800 68.000 ;
        RECT 110.200 67.900 110.600 69.900 ;
        RECT 112.600 67.900 113.000 69.900 ;
        RECT 113.300 68.200 113.700 68.600 ;
        RECT 104.700 67.200 105.000 67.900 ;
        RECT 105.500 67.700 107.300 67.900 ;
        RECT 107.900 67.700 109.700 67.900 ;
        RECT 106.600 67.200 107.000 67.400 ;
        RECT 108.200 67.200 108.600 67.400 ;
        RECT 110.200 67.200 110.500 67.900 ;
        RECT 104.600 66.800 105.900 67.200 ;
        RECT 106.600 67.100 107.400 67.200 ;
        RECT 107.800 67.100 108.600 67.200 ;
        RECT 106.600 66.900 108.600 67.100 ;
        RECT 107.000 66.800 108.200 66.900 ;
        RECT 109.300 66.800 110.600 67.200 ;
        RECT 111.000 67.100 111.400 67.200 ;
        RECT 111.800 67.100 112.200 67.200 ;
        RECT 111.000 66.800 112.200 67.100 ;
        RECT 104.600 66.100 105.000 66.200 ;
        RECT 100.600 65.800 105.000 66.100 ;
        RECT 100.600 65.200 100.900 65.800 ;
        RECT 100.600 65.100 101.000 65.200 ;
        RECT 89.400 64.800 90.500 65.100 ;
        RECT 89.400 61.100 89.800 64.800 ;
        RECT 92.300 61.100 93.300 65.100 ;
        RECT 95.000 64.800 95.700 65.100 ;
        RECT 96.000 64.800 96.500 65.100 ;
        RECT 95.400 64.200 95.700 64.800 ;
        RECT 95.400 63.800 95.800 64.200 ;
        RECT 96.100 61.100 96.500 64.800 ;
        RECT 99.500 64.800 100.000 65.100 ;
        RECT 100.300 64.800 101.000 65.100 ;
        RECT 99.500 62.200 99.900 64.800 ;
        RECT 100.300 64.200 100.600 64.800 ;
        RECT 100.200 63.800 100.600 64.200 ;
        RECT 99.000 61.800 99.900 62.200 ;
        RECT 99.500 61.100 99.900 61.800 ;
        RECT 103.800 61.100 104.200 65.800 ;
        RECT 104.600 65.100 105.000 65.200 ;
        RECT 105.600 65.100 105.900 66.800 ;
        RECT 106.200 66.100 106.600 66.600 ;
        RECT 108.600 66.100 109.000 66.600 ;
        RECT 106.200 65.800 109.000 66.100 ;
        RECT 109.300 65.100 109.600 66.800 ;
        RECT 111.800 66.400 112.200 66.800 ;
        RECT 110.200 66.100 110.600 66.200 ;
        RECT 111.000 66.100 111.400 66.200 ;
        RECT 112.600 66.100 112.900 67.900 ;
        RECT 113.400 67.800 113.800 68.200 ;
        RECT 116.000 67.100 116.400 69.900 ;
        RECT 118.000 67.100 118.400 69.900 ;
        RECT 116.000 66.900 116.900 67.100 ;
        RECT 116.100 66.800 116.900 66.900 ;
        RECT 113.400 66.100 113.800 66.200 ;
        RECT 110.200 65.800 111.800 66.100 ;
        RECT 112.600 65.800 113.800 66.100 ;
        RECT 115.000 65.800 115.800 66.200 ;
        RECT 111.400 65.600 111.800 65.800 ;
        RECT 110.200 65.100 110.600 65.200 ;
        RECT 113.400 65.100 113.700 65.800 ;
        RECT 104.600 64.800 105.300 65.100 ;
        RECT 105.600 64.800 106.100 65.100 ;
        RECT 105.000 64.200 105.300 64.800 ;
        RECT 105.000 63.800 105.400 64.200 ;
        RECT 105.700 62.200 106.100 64.800 ;
        RECT 109.100 64.800 109.600 65.100 ;
        RECT 109.900 64.800 110.600 65.100 ;
        RECT 111.000 64.800 113.000 65.100 ;
        RECT 109.100 62.200 109.500 64.800 ;
        RECT 109.900 64.200 110.200 64.800 ;
        RECT 109.800 63.800 110.200 64.200 ;
        RECT 105.700 61.800 106.600 62.200 ;
        RECT 108.600 61.800 109.500 62.200 ;
        RECT 105.700 61.100 106.100 61.800 ;
        RECT 109.100 61.100 109.500 61.800 ;
        RECT 111.000 61.100 111.400 64.800 ;
        RECT 112.600 61.100 113.000 64.800 ;
        RECT 113.400 61.100 113.800 65.100 ;
        RECT 114.200 64.800 114.600 65.600 ;
        RECT 116.600 65.200 116.900 66.800 ;
        RECT 117.500 66.900 118.400 67.100 ;
        RECT 122.400 67.100 122.800 69.900 ;
        RECT 125.400 67.800 125.800 69.900 ;
        RECT 126.100 68.200 126.500 68.600 ;
        RECT 126.200 67.800 126.600 68.200 ;
        RECT 122.400 66.900 123.300 67.100 ;
        RECT 117.500 66.800 118.300 66.900 ;
        RECT 122.500 66.800 123.300 66.900 ;
        RECT 117.500 65.200 117.800 66.800 ;
        RECT 118.600 65.800 119.400 66.200 ;
        RECT 121.400 65.800 122.200 66.200 ;
        RECT 116.600 64.800 117.000 65.200 ;
        RECT 117.400 64.800 117.800 65.200 ;
        RECT 115.800 63.800 116.200 64.600 ;
        RECT 116.600 63.500 116.900 64.800 ;
        RECT 115.100 63.200 116.900 63.500 ;
        RECT 115.100 63.100 115.400 63.200 ;
        RECT 115.000 61.100 115.400 63.100 ;
        RECT 116.600 63.100 116.900 63.200 ;
        RECT 117.500 63.500 117.800 64.800 ;
        RECT 118.200 64.100 118.600 65.200 ;
        RECT 119.800 64.800 120.200 65.600 ;
        RECT 120.600 64.800 121.000 65.600 ;
        RECT 123.000 65.200 123.300 66.800 ;
        RECT 124.600 66.400 125.000 67.200 ;
        RECT 123.800 66.100 124.200 66.200 ;
        RECT 125.400 66.100 125.700 67.800 ;
        RECT 128.800 67.100 129.200 69.900 ;
        RECT 132.000 67.100 132.400 69.900 ;
        RECT 135.200 67.100 135.600 69.900 ;
        RECT 138.200 67.900 138.600 69.900 ;
        RECT 138.900 68.200 139.300 68.600 ;
        RECT 128.800 66.900 129.700 67.100 ;
        RECT 132.000 66.900 132.900 67.100 ;
        RECT 135.200 66.900 136.100 67.100 ;
        RECT 128.900 66.800 129.700 66.900 ;
        RECT 132.100 66.800 132.900 66.900 ;
        RECT 135.300 66.800 136.100 66.900 ;
        RECT 126.200 66.100 126.600 66.200 ;
        RECT 123.800 65.800 124.600 66.100 ;
        RECT 125.400 65.800 126.600 66.100 ;
        RECT 127.800 65.800 128.600 66.200 ;
        RECT 124.200 65.600 124.600 65.800 ;
        RECT 123.000 64.800 123.400 65.200 ;
        RECT 126.200 65.100 126.500 65.800 ;
        RECT 123.800 64.800 125.800 65.100 ;
        RECT 118.200 63.800 121.700 64.100 ;
        RECT 122.200 63.800 122.600 64.600 ;
        RECT 121.400 63.500 121.700 63.800 ;
        RECT 123.000 63.500 123.300 64.800 ;
        RECT 117.500 63.200 119.300 63.500 ;
        RECT 117.500 63.100 117.800 63.200 ;
        RECT 116.600 61.100 117.000 63.100 ;
        RECT 117.400 61.100 117.800 63.100 ;
        RECT 119.000 63.100 119.300 63.200 ;
        RECT 121.400 63.200 123.300 63.500 ;
        RECT 119.000 61.100 119.400 63.100 ;
        RECT 121.400 61.100 121.800 63.200 ;
        RECT 123.000 63.100 123.300 63.200 ;
        RECT 123.000 61.100 123.400 63.100 ;
        RECT 123.800 61.100 124.200 64.800 ;
        RECT 125.400 61.100 125.800 64.800 ;
        RECT 126.200 61.100 126.600 65.100 ;
        RECT 127.000 64.800 127.400 65.600 ;
        RECT 129.400 65.200 129.700 66.800 ;
        RECT 131.000 65.800 131.800 66.200 ;
        RECT 129.400 64.800 129.800 65.200 ;
        RECT 130.200 64.800 130.600 65.600 ;
        RECT 132.600 65.200 132.900 66.800 ;
        RECT 134.200 65.800 135.000 66.200 ;
        RECT 131.000 65.100 131.400 65.200 ;
        RECT 131.000 64.800 132.200 65.100 ;
        RECT 128.600 63.800 129.000 64.600 ;
        RECT 129.400 64.100 129.700 64.800 ;
        RECT 131.800 64.100 132.200 64.800 ;
        RECT 129.400 63.800 132.200 64.100 ;
        RECT 132.600 64.800 133.000 65.200 ;
        RECT 133.400 64.800 133.800 65.600 ;
        RECT 135.800 65.200 136.100 66.800 ;
        RECT 137.400 66.400 137.800 67.200 ;
        RECT 136.600 66.100 137.000 66.200 ;
        RECT 138.200 66.100 138.500 67.900 ;
        RECT 139.000 67.800 139.400 68.200 ;
        RECT 140.400 67.100 140.800 69.900 ;
        RECT 143.600 67.100 144.000 69.900 ;
        RECT 146.200 67.900 146.600 69.900 ;
        RECT 148.400 69.200 149.200 69.900 ;
        RECT 147.800 68.800 149.200 69.200 ;
        RECT 148.400 68.100 149.200 68.800 ;
        RECT 146.200 67.600 147.400 67.900 ;
        RECT 147.000 67.500 147.400 67.600 ;
        RECT 147.700 67.400 148.100 67.800 ;
        RECT 147.700 67.200 148.000 67.400 ;
        RECT 139.900 66.900 140.800 67.100 ;
        RECT 143.100 66.900 144.000 67.100 ;
        RECT 139.900 66.800 140.700 66.900 ;
        RECT 143.100 66.800 143.900 66.900 ;
        RECT 146.200 66.800 147.000 67.200 ;
        RECT 147.600 66.800 148.000 67.200 ;
        RECT 148.400 67.100 148.700 68.100 ;
        RECT 151.000 67.900 151.400 69.900 ;
        RECT 149.000 67.400 149.800 67.800 ;
        RECT 150.100 67.600 151.400 67.900 ;
        RECT 150.100 67.500 150.500 67.600 ;
        RECT 150.600 67.100 151.400 67.200 ;
        RECT 148.400 66.800 148.900 67.100 ;
        RECT 150.300 67.000 151.400 67.100 ;
        RECT 139.000 66.100 139.400 66.200 ;
        RECT 136.600 65.800 137.400 66.100 ;
        RECT 138.200 65.800 139.400 66.100 ;
        RECT 137.000 65.600 137.400 65.800 ;
        RECT 135.800 64.800 136.200 65.200 ;
        RECT 139.000 65.100 139.300 65.800 ;
        RECT 139.900 65.200 140.200 66.800 ;
        RECT 141.000 65.800 141.800 66.200 ;
        RECT 136.600 64.800 138.600 65.100 ;
        RECT 129.400 63.500 129.700 63.800 ;
        RECT 132.600 63.500 132.900 64.800 ;
        RECT 135.000 63.800 135.400 64.600 ;
        RECT 135.800 63.500 136.100 64.800 ;
        RECT 127.900 63.200 129.700 63.500 ;
        RECT 127.900 63.100 128.200 63.200 ;
        RECT 127.800 61.100 128.200 63.100 ;
        RECT 129.400 63.100 129.700 63.200 ;
        RECT 131.100 63.200 132.900 63.500 ;
        RECT 131.100 63.100 131.400 63.200 ;
        RECT 129.400 61.100 129.800 63.100 ;
        RECT 131.000 61.100 131.400 63.100 ;
        RECT 132.600 63.100 132.900 63.200 ;
        RECT 134.300 63.200 136.100 63.500 ;
        RECT 134.300 63.100 134.600 63.200 ;
        RECT 132.600 61.100 133.000 63.100 ;
        RECT 134.200 61.100 134.600 63.100 ;
        RECT 135.800 63.100 136.100 63.200 ;
        RECT 135.800 61.100 136.200 63.100 ;
        RECT 136.600 61.100 137.000 64.800 ;
        RECT 138.200 61.100 138.600 64.800 ;
        RECT 139.000 61.100 139.400 65.100 ;
        RECT 139.800 64.800 140.200 65.200 ;
        RECT 142.200 64.800 142.600 65.600 ;
        RECT 143.100 65.200 143.400 66.800 ;
        RECT 148.600 66.200 148.900 66.800 ;
        RECT 149.200 66.800 151.400 67.000 ;
        RECT 149.200 66.700 150.600 66.800 ;
        RECT 149.200 66.600 149.600 66.700 ;
        RECT 144.200 65.800 145.000 66.200 ;
        RECT 148.600 65.800 149.000 66.200 ;
        RECT 149.900 66.100 150.300 66.200 ;
        RECT 149.500 65.800 150.300 66.100 ;
        RECT 143.000 64.800 143.400 65.200 ;
        RECT 145.400 64.800 145.800 65.600 ;
        RECT 148.600 65.100 148.900 65.800 ;
        RECT 149.500 65.700 149.900 65.800 ;
        RECT 146.200 64.800 147.400 65.100 ;
        RECT 139.900 63.500 140.200 64.800 ;
        RECT 140.600 63.800 141.000 64.600 ;
        RECT 143.100 63.500 143.400 64.800 ;
        RECT 143.800 63.800 144.200 64.600 ;
        RECT 139.900 63.200 141.700 63.500 ;
        RECT 139.900 63.100 140.200 63.200 ;
        RECT 139.800 61.100 140.200 63.100 ;
        RECT 141.400 63.100 141.700 63.200 ;
        RECT 143.100 63.200 144.900 63.500 ;
        RECT 143.100 63.100 143.400 63.200 ;
        RECT 141.400 61.100 141.800 63.100 ;
        RECT 143.000 61.100 143.400 63.100 ;
        RECT 144.600 63.100 144.900 63.200 ;
        RECT 144.600 61.100 145.000 63.100 ;
        RECT 146.200 61.100 146.600 64.800 ;
        RECT 147.000 64.700 147.400 64.800 ;
        RECT 148.400 62.200 149.200 65.100 ;
        RECT 150.100 64.800 151.400 65.100 ;
        RECT 150.100 64.700 150.500 64.800 ;
        RECT 148.400 61.800 149.800 62.200 ;
        RECT 148.400 61.100 149.200 61.800 ;
        RECT 151.000 61.100 151.400 64.800 ;
        RECT 0.600 56.200 1.000 59.900 ;
        RECT 1.300 56.200 1.700 56.300 ;
        RECT 0.600 55.900 1.700 56.200 ;
        RECT 2.800 56.200 3.600 59.900 ;
        RECT 4.600 56.200 5.000 56.300 ;
        RECT 5.400 56.200 5.800 59.900 ;
        RECT 2.800 55.900 3.800 56.200 ;
        RECT 4.600 55.900 5.800 56.200 ;
        RECT 1.400 55.600 1.700 55.900 ;
        RECT 1.400 55.300 3.100 55.600 ;
        RECT 2.700 55.200 3.100 55.300 ;
        RECT 3.500 55.200 3.800 55.900 ;
        RECT 6.200 55.700 6.600 59.900 ;
        RECT 8.400 58.200 8.800 59.900 ;
        RECT 7.800 57.900 8.800 58.200 ;
        RECT 10.600 57.900 11.000 59.900 ;
        RECT 12.700 57.900 13.300 59.900 ;
        RECT 7.800 57.500 8.200 57.900 ;
        RECT 10.600 57.600 10.900 57.900 ;
        RECT 9.500 57.300 11.300 57.600 ;
        RECT 12.600 57.500 13.000 57.900 ;
        RECT 9.500 57.200 9.900 57.300 ;
        RECT 10.900 57.200 11.300 57.300 ;
        RECT 7.800 56.500 8.200 56.600 ;
        RECT 10.100 56.500 10.500 56.600 ;
        RECT 7.800 56.200 10.500 56.500 ;
        RECT 10.800 56.500 11.900 56.800 ;
        RECT 10.800 55.900 11.100 56.500 ;
        RECT 11.500 56.400 11.900 56.500 ;
        RECT 12.700 56.600 13.400 57.000 ;
        RECT 12.700 56.100 13.000 56.600 ;
        RECT 8.700 55.700 11.100 55.900 ;
        RECT 6.200 55.600 11.100 55.700 ;
        RECT 11.800 55.800 13.000 56.100 ;
        RECT 6.200 55.500 9.100 55.600 ;
        RECT 6.200 55.400 9.000 55.500 ;
        RECT 11.800 55.200 12.100 55.800 ;
        RECT 15.000 55.600 15.400 59.900 ;
        RECT 15.800 56.200 16.200 59.900 ;
        RECT 18.000 59.200 18.800 59.900 ;
        RECT 18.000 58.800 19.400 59.200 ;
        RECT 16.500 56.200 16.900 56.300 ;
        RECT 15.800 55.900 16.900 56.200 ;
        RECT 18.000 56.200 18.800 58.800 ;
        RECT 19.800 56.200 20.200 56.300 ;
        RECT 20.600 56.200 21.000 59.900 ;
        RECT 18.000 55.900 19.000 56.200 ;
        RECT 19.800 55.900 21.000 56.200 ;
        RECT 13.300 55.300 15.400 55.600 ;
        RECT 16.600 55.600 16.900 55.900 ;
        RECT 16.600 55.300 18.300 55.600 ;
        RECT 13.300 55.200 13.700 55.300 ;
        RECT 1.600 54.900 2.000 55.000 ;
        RECT 3.500 54.900 4.200 55.200 ;
        RECT 9.400 55.100 9.800 55.200 ;
        RECT 1.600 54.600 2.900 54.900 ;
        RECT 2.600 54.300 2.900 54.600 ;
        RECT 3.300 54.800 4.200 54.900 ;
        RECT 7.300 54.800 9.800 55.100 ;
        RECT 11.800 54.800 12.200 55.200 ;
        RECT 14.100 54.900 14.500 55.000 ;
        RECT 3.300 54.600 3.800 54.800 ;
        RECT 7.300 54.700 7.700 54.800 ;
        RECT 8.600 54.700 9.000 54.800 ;
        RECT 0.600 54.100 1.400 54.200 ;
        RECT 0.600 53.800 2.300 54.100 ;
        RECT 2.600 53.900 3.000 54.300 ;
        RECT 2.000 53.600 2.300 53.800 ;
        RECT 1.300 53.400 1.700 53.500 ;
        RECT 0.600 53.100 1.700 53.400 ;
        RECT 2.000 53.300 3.000 53.600 ;
        RECT 2.200 53.200 3.000 53.300 ;
        RECT 0.600 51.100 1.000 53.100 ;
        RECT 3.300 52.900 3.600 54.600 ;
        RECT 8.100 54.200 8.500 54.300 ;
        RECT 11.800 54.200 12.100 54.800 ;
        RECT 12.600 54.600 14.500 54.900 ;
        RECT 12.600 54.500 13.000 54.600 ;
        RECT 4.000 53.800 4.400 54.200 ;
        RECT 5.000 53.800 5.800 54.200 ;
        RECT 6.600 53.900 12.100 54.200 ;
        RECT 6.600 53.800 7.400 53.900 ;
        RECT 4.000 53.600 4.300 53.800 ;
        RECT 3.900 53.200 4.300 53.600 ;
        RECT 4.600 53.400 5.000 53.500 ;
        RECT 4.600 53.100 5.800 53.400 ;
        RECT 2.800 51.100 3.600 52.900 ;
        RECT 5.400 51.100 5.800 53.100 ;
        RECT 6.200 51.100 6.600 53.500 ;
        RECT 8.700 52.800 9.000 53.900 ;
        RECT 11.500 53.800 11.900 53.900 ;
        RECT 15.000 53.600 15.400 55.300 ;
        RECT 17.900 55.200 18.300 55.300 ;
        RECT 18.700 55.200 19.000 55.900 ;
        RECT 16.800 54.900 17.200 55.000 ;
        RECT 18.700 54.900 19.400 55.200 ;
        RECT 16.800 54.600 18.100 54.900 ;
        RECT 17.800 54.300 18.100 54.600 ;
        RECT 18.500 54.800 19.400 54.900 ;
        RECT 18.500 54.600 19.000 54.800 ;
        RECT 15.800 54.100 16.600 54.200 ;
        RECT 15.800 53.800 17.500 54.100 ;
        RECT 17.800 53.900 18.200 54.300 ;
        RECT 13.500 53.300 15.400 53.600 ;
        RECT 17.200 53.600 17.500 53.800 ;
        RECT 16.500 53.400 16.900 53.500 ;
        RECT 13.500 53.200 13.900 53.300 ;
        RECT 7.800 52.100 8.200 52.500 ;
        RECT 8.600 52.400 9.000 52.800 ;
        RECT 9.500 52.700 9.900 52.800 ;
        RECT 9.500 52.400 10.900 52.700 ;
        RECT 10.600 52.100 10.900 52.400 ;
        RECT 12.600 52.100 13.000 52.500 ;
        RECT 7.800 51.800 8.800 52.100 ;
        RECT 8.400 51.100 8.800 51.800 ;
        RECT 10.600 51.100 11.000 52.100 ;
        RECT 12.600 51.800 13.300 52.100 ;
        RECT 12.700 51.100 13.300 51.800 ;
        RECT 15.000 51.100 15.400 53.300 ;
        RECT 15.800 53.100 16.900 53.400 ;
        RECT 17.200 53.300 18.200 53.600 ;
        RECT 17.400 53.200 18.200 53.300 ;
        RECT 15.800 51.100 16.200 53.100 ;
        RECT 18.500 52.900 18.800 54.600 ;
        RECT 19.200 53.800 19.600 54.200 ;
        RECT 20.200 53.800 21.000 54.200 ;
        RECT 19.200 53.600 19.500 53.800 ;
        RECT 19.100 53.200 19.500 53.600 ;
        RECT 19.800 53.400 20.200 53.500 ;
        RECT 21.400 53.400 21.800 54.200 ;
        RECT 19.800 53.100 21.000 53.400 ;
        RECT 18.000 51.100 18.800 52.900 ;
        RECT 20.600 51.100 21.000 53.100 ;
        RECT 22.200 53.100 22.600 59.900 ;
        RECT 23.000 56.100 23.400 56.600 ;
        RECT 23.800 56.100 24.200 56.200 ;
        RECT 23.000 55.800 24.200 56.100 ;
        RECT 23.800 53.100 24.200 53.200 ;
        RECT 22.200 52.800 24.200 53.100 ;
        RECT 22.700 51.100 23.100 52.800 ;
        RECT 23.800 52.400 24.200 52.800 ;
        RECT 24.600 51.100 25.000 59.900 ;
        RECT 26.700 56.300 27.100 59.900 ;
        RECT 29.100 56.300 29.500 59.900 ;
        RECT 26.200 55.900 27.100 56.300 ;
        RECT 28.600 55.900 29.500 56.300 ;
        RECT 26.300 54.200 26.600 55.900 ;
        RECT 27.000 54.800 27.400 55.600 ;
        RECT 28.700 54.200 29.000 55.900 ;
        RECT 29.400 54.800 29.800 55.600 ;
        RECT 26.200 53.800 26.600 54.200 ;
        RECT 28.600 53.800 29.000 54.200 ;
        RECT 25.400 52.400 25.800 53.200 ;
        RECT 26.300 53.100 26.600 53.800 ;
        RECT 27.800 53.100 28.200 53.200 ;
        RECT 28.700 53.100 29.000 53.800 ;
        RECT 30.200 53.100 30.600 53.200 ;
        RECT 26.200 52.800 28.200 53.100 ;
        RECT 28.600 52.800 30.600 53.100 ;
        RECT 26.300 52.100 26.600 52.800 ;
        RECT 27.800 52.400 28.200 52.800 ;
        RECT 28.700 52.100 29.000 52.800 ;
        RECT 30.200 52.400 30.600 52.800 ;
        RECT 26.200 51.100 26.600 52.100 ;
        RECT 28.600 51.100 29.000 52.100 ;
        RECT 31.000 51.100 31.400 59.900 ;
        RECT 32.600 55.600 33.000 59.900 ;
        RECT 34.200 55.600 34.600 59.900 ;
        RECT 35.800 55.600 36.200 59.900 ;
        RECT 37.400 55.600 37.800 59.900 ;
        RECT 31.800 55.200 33.000 55.600 ;
        RECT 31.800 53.800 32.200 55.200 ;
        RECT 32.600 54.800 33.000 55.200 ;
        RECT 33.500 55.200 34.600 55.600 ;
        RECT 35.100 55.200 36.200 55.600 ;
        RECT 36.900 55.200 37.800 55.600 ;
        RECT 39.000 55.700 39.400 59.900 ;
        RECT 41.200 58.200 41.600 59.900 ;
        RECT 40.600 57.900 41.600 58.200 ;
        RECT 43.400 57.900 43.800 59.900 ;
        RECT 45.500 57.900 46.100 59.900 ;
        RECT 40.600 57.500 41.000 57.900 ;
        RECT 43.400 57.600 43.700 57.900 ;
        RECT 42.300 57.300 44.100 57.600 ;
        RECT 45.400 57.500 45.800 57.900 ;
        RECT 42.300 57.200 42.700 57.300 ;
        RECT 43.700 57.200 44.100 57.300 ;
        RECT 40.600 56.500 41.000 56.600 ;
        RECT 42.900 56.500 43.300 56.600 ;
        RECT 40.600 56.200 43.300 56.500 ;
        RECT 43.600 56.500 44.700 56.800 ;
        RECT 43.600 55.900 43.900 56.500 ;
        RECT 44.300 56.400 44.700 56.500 ;
        RECT 45.500 56.600 46.200 57.000 ;
        RECT 45.500 56.100 45.800 56.600 ;
        RECT 41.500 55.700 43.900 55.900 ;
        RECT 39.000 55.600 43.900 55.700 ;
        RECT 44.600 55.800 45.800 56.100 ;
        RECT 39.000 55.500 41.900 55.600 ;
        RECT 39.000 55.400 41.800 55.500 ;
        RECT 33.500 54.500 33.900 55.200 ;
        RECT 35.100 54.500 35.500 55.200 ;
        RECT 36.900 54.500 37.300 55.200 ;
        RECT 42.200 55.100 42.600 55.200 ;
        RECT 40.100 54.800 42.600 55.100 ;
        RECT 40.100 54.700 40.500 54.800 ;
        RECT 32.600 54.100 33.900 54.500 ;
        RECT 34.300 54.100 35.500 54.500 ;
        RECT 36.000 54.100 37.300 54.500 ;
        RECT 40.900 54.200 41.300 54.300 ;
        RECT 44.600 54.200 44.900 55.800 ;
        RECT 47.800 55.600 48.200 59.900 ;
        RECT 50.200 56.200 50.600 59.900 ;
        RECT 51.800 56.200 52.200 59.900 ;
        RECT 50.200 55.900 52.200 56.200 ;
        RECT 52.600 55.900 53.000 59.900 ;
        RECT 53.400 57.900 53.800 59.900 ;
        RECT 53.500 57.800 53.800 57.900 ;
        RECT 55.000 57.900 55.400 59.900 ;
        RECT 55.000 57.800 55.300 57.900 ;
        RECT 53.500 57.500 55.300 57.800 ;
        RECT 53.500 56.200 53.800 57.500 ;
        RECT 46.100 55.300 48.200 55.600 ;
        RECT 46.100 55.200 46.500 55.300 ;
        RECT 46.900 54.900 47.300 55.000 ;
        RECT 45.400 54.600 47.300 54.900 ;
        RECT 45.400 54.500 45.800 54.600 ;
        RECT 33.500 53.800 33.900 54.100 ;
        RECT 35.100 53.800 35.500 54.100 ;
        RECT 36.900 53.800 37.300 54.100 ;
        RECT 39.400 53.900 44.900 54.200 ;
        RECT 47.800 54.100 48.200 55.300 ;
        RECT 50.600 55.200 51.000 55.400 ;
        RECT 52.600 55.200 52.900 55.900 ;
        RECT 53.400 55.800 53.800 56.200 ;
        RECT 54.200 57.100 54.600 57.200 ;
        RECT 57.400 57.100 57.800 59.900 ;
        RECT 54.200 56.800 57.800 57.100 ;
        RECT 54.200 56.100 54.600 56.800 ;
        RECT 55.000 56.100 55.400 56.200 ;
        RECT 54.200 55.800 55.400 56.100 ;
        RECT 50.200 54.900 51.000 55.200 ;
        RECT 51.800 54.900 53.000 55.200 ;
        RECT 50.200 54.800 50.600 54.900 ;
        RECT 51.000 54.100 51.400 54.600 ;
        RECT 39.400 53.800 40.200 53.900 ;
        RECT 31.800 53.400 33.000 53.800 ;
        RECT 33.500 53.400 34.600 53.800 ;
        RECT 35.100 53.400 36.200 53.800 ;
        RECT 36.900 53.400 37.800 53.800 ;
        RECT 32.600 51.100 33.000 53.400 ;
        RECT 34.200 51.100 34.600 53.400 ;
        RECT 35.800 51.100 36.200 53.400 ;
        RECT 37.400 51.100 37.800 53.400 ;
        RECT 39.000 51.100 39.400 53.500 ;
        RECT 41.500 52.800 41.800 53.900 ;
        RECT 43.000 53.800 43.400 53.900 ;
        RECT 44.300 53.800 44.700 53.900 ;
        RECT 47.800 53.800 51.400 54.100 ;
        RECT 47.800 53.600 48.200 53.800 ;
        RECT 46.300 53.300 48.200 53.600 ;
        RECT 46.300 53.200 46.700 53.300 ;
        RECT 40.600 52.100 41.000 52.500 ;
        RECT 41.400 52.400 41.800 52.800 ;
        RECT 42.300 52.700 42.700 52.800 ;
        RECT 42.300 52.400 43.700 52.700 ;
        RECT 43.400 52.100 43.700 52.400 ;
        RECT 45.400 52.100 45.800 52.500 ;
        RECT 40.600 51.800 41.600 52.100 ;
        RECT 41.200 51.100 41.600 51.800 ;
        RECT 43.400 51.100 43.800 52.100 ;
        RECT 45.400 51.800 46.100 52.100 ;
        RECT 45.500 51.100 46.100 51.800 ;
        RECT 47.800 51.100 48.200 53.300 ;
        RECT 51.800 53.100 52.100 54.900 ;
        RECT 52.600 54.800 53.000 54.900 ;
        RECT 53.500 54.200 53.800 55.800 ;
        RECT 55.800 55.400 56.200 56.200 ;
        RECT 54.600 54.800 55.400 55.200 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 56.600 54.200 56.900 54.800 ;
        RECT 53.500 54.100 54.300 54.200 ;
        RECT 53.500 53.900 54.400 54.100 ;
        RECT 51.800 51.100 52.200 53.100 ;
        RECT 52.600 52.800 53.000 53.200 ;
        RECT 52.500 52.400 52.900 52.800 ;
        RECT 54.000 51.100 54.400 53.900 ;
        RECT 56.600 53.400 57.000 54.200 ;
        RECT 57.400 53.100 57.800 56.800 ;
        RECT 58.200 55.800 58.600 56.600 ;
        RECT 59.000 53.400 59.400 54.200 ;
        RECT 59.800 53.100 60.200 59.900 ;
        RECT 60.600 55.800 61.000 56.600 ;
        RECT 61.400 53.400 61.800 54.200 ;
        RECT 62.200 53.100 62.600 59.900 ;
        RECT 63.000 55.800 63.400 56.600 ;
        RECT 63.800 55.800 64.200 56.600 ;
        RECT 64.600 53.100 65.000 59.900 ;
        RECT 66.200 56.200 66.600 59.900 ;
        RECT 67.800 56.400 68.200 59.900 ;
        RECT 70.700 59.200 71.100 59.900 ;
        RECT 70.200 58.800 71.100 59.200 ;
        RECT 66.200 55.900 67.500 56.200 ;
        RECT 67.800 55.900 68.300 56.400 ;
        RECT 70.700 56.200 71.100 58.800 ;
        RECT 71.400 56.800 71.800 57.200 ;
        RECT 71.500 56.200 71.800 56.800 ;
        RECT 70.700 55.900 71.200 56.200 ;
        RECT 71.500 55.900 72.200 56.200 ;
        RECT 65.400 54.800 65.800 55.200 ;
        RECT 66.200 54.800 66.700 55.200 ;
        RECT 65.400 54.200 65.700 54.800 ;
        RECT 66.300 54.400 66.700 54.800 ;
        RECT 67.200 54.900 67.500 55.900 ;
        RECT 67.200 54.500 67.700 54.900 ;
        RECT 65.400 53.400 65.800 54.200 ;
        RECT 67.200 53.700 67.500 54.500 ;
        RECT 68.000 54.200 68.300 55.900 ;
        RECT 70.200 54.400 70.600 55.200 ;
        RECT 70.900 54.200 71.200 55.900 ;
        RECT 71.800 55.800 72.200 55.900 ;
        RECT 67.800 54.100 68.300 54.200 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 67.800 53.800 69.000 54.100 ;
        RECT 69.400 54.100 69.800 54.200 ;
        RECT 69.400 53.800 70.200 54.100 ;
        RECT 70.900 53.800 72.200 54.200 ;
        RECT 66.200 53.400 67.500 53.700 ;
        RECT 57.400 52.800 58.300 53.100 ;
        RECT 59.800 52.800 60.700 53.100 ;
        RECT 62.200 52.800 63.100 53.100 ;
        RECT 57.900 52.200 58.300 52.800 ;
        RECT 60.300 52.200 60.700 52.800 ;
        RECT 62.700 52.200 63.100 52.800 ;
        RECT 64.100 52.800 65.000 53.100 ;
        RECT 64.100 52.200 64.500 52.800 ;
        RECT 57.900 51.800 58.600 52.200 ;
        RECT 60.300 51.800 61.000 52.200 ;
        RECT 62.700 51.800 63.400 52.200 ;
        RECT 64.100 51.800 65.000 52.200 ;
        RECT 57.900 51.100 58.300 51.800 ;
        RECT 60.300 51.100 60.700 51.800 ;
        RECT 62.700 51.100 63.100 51.800 ;
        RECT 64.100 51.100 64.500 51.800 ;
        RECT 66.200 51.100 66.600 53.400 ;
        RECT 68.000 53.100 68.300 53.800 ;
        RECT 69.800 53.600 70.200 53.800 ;
        RECT 69.500 53.100 71.300 53.300 ;
        RECT 71.800 53.100 72.100 53.800 ;
        RECT 72.600 53.400 73.000 54.200 ;
        RECT 73.400 54.100 73.800 59.900 ;
        RECT 74.200 56.100 74.600 56.600 ;
        RECT 75.000 56.100 75.400 56.600 ;
        RECT 74.200 55.800 75.400 56.100 ;
        RECT 74.200 55.200 74.500 55.800 ;
        RECT 74.200 54.800 74.600 55.200 ;
        RECT 74.200 54.100 74.600 54.200 ;
        RECT 73.400 53.800 74.600 54.100 ;
        RECT 73.400 53.100 73.800 53.800 ;
        RECT 75.800 53.100 76.200 59.900 ;
        RECT 76.600 53.400 77.000 54.200 ;
        RECT 77.400 53.400 77.800 54.200 ;
        RECT 67.800 52.800 68.300 53.100 ;
        RECT 69.400 53.000 71.400 53.100 ;
        RECT 67.800 51.100 68.200 52.800 ;
        RECT 69.400 51.100 69.800 53.000 ;
        RECT 71.000 51.100 71.400 53.000 ;
        RECT 71.800 51.100 72.200 53.100 ;
        RECT 73.400 52.800 74.300 53.100 ;
        RECT 73.900 51.100 74.300 52.800 ;
        RECT 75.300 52.800 76.200 53.100 ;
        RECT 78.200 53.100 78.600 59.900 ;
        RECT 79.000 56.100 79.400 56.600 ;
        RECT 79.800 56.100 80.200 57.200 ;
        RECT 79.000 55.800 80.200 56.100 ;
        RECT 80.600 53.100 81.000 59.900 ;
        RECT 83.500 56.300 83.900 59.900 ;
        RECT 83.000 55.900 83.900 56.300 ;
        RECT 85.900 55.900 86.900 59.900 ;
        RECT 88.600 55.900 89.000 59.900 ;
        RECT 89.400 56.200 89.800 59.900 ;
        RECT 91.000 56.200 91.400 59.900 ;
        RECT 92.600 57.900 93.000 59.900 ;
        RECT 92.700 57.800 93.000 57.900 ;
        RECT 94.200 57.900 94.600 59.900 ;
        RECT 95.000 57.900 95.400 59.900 ;
        RECT 94.200 57.800 94.500 57.900 ;
        RECT 92.700 57.500 94.500 57.800 ;
        RECT 93.400 56.400 93.800 57.200 ;
        RECT 94.200 56.200 94.500 57.500 ;
        RECT 95.100 57.800 95.400 57.900 ;
        RECT 96.600 57.900 97.000 59.900 ;
        RECT 96.600 57.800 96.900 57.900 ;
        RECT 95.100 57.500 96.900 57.800 ;
        RECT 95.100 56.200 95.400 57.500 ;
        RECT 95.800 56.400 96.200 57.200 ;
        RECT 98.200 56.200 98.600 59.900 ;
        RECT 99.800 56.200 100.200 59.900 ;
        RECT 89.400 55.900 91.400 56.200 ;
        RECT 83.100 54.200 83.400 55.900 ;
        RECT 83.800 54.800 84.200 55.600 ;
        RECT 84.600 55.100 85.000 55.200 ;
        RECT 85.400 55.100 85.800 55.200 ;
        RECT 84.600 54.800 85.800 55.100 ;
        RECT 85.400 54.400 85.800 54.800 ;
        RECT 86.200 54.200 86.500 55.900 ;
        RECT 88.700 55.200 89.000 55.900 ;
        RECT 91.800 55.400 92.200 56.200 ;
        RECT 94.200 55.800 94.600 56.200 ;
        RECT 95.000 55.800 95.400 56.200 ;
        RECT 90.600 55.200 91.000 55.400 ;
        RECT 87.000 54.400 87.400 55.200 ;
        RECT 88.600 54.900 89.800 55.200 ;
        RECT 90.600 54.900 91.400 55.200 ;
        RECT 88.600 54.800 89.000 54.900 ;
        RECT 81.400 54.100 81.800 54.200 ;
        RECT 82.200 54.100 82.600 54.200 ;
        RECT 81.400 53.800 82.600 54.100 ;
        RECT 83.000 53.800 83.400 54.200 ;
        RECT 83.800 54.100 84.200 54.200 ;
        RECT 84.600 54.100 85.000 54.200 ;
        RECT 86.200 54.100 86.600 54.200 ;
        RECT 83.800 53.800 85.400 54.100 ;
        RECT 86.200 53.800 87.400 54.100 ;
        RECT 87.800 53.800 88.200 54.600 ;
        RECT 81.400 53.400 81.800 53.800 ;
        RECT 78.200 52.800 79.100 53.100 ;
        RECT 75.300 52.200 75.700 52.800 ;
        RECT 78.700 52.200 79.100 52.800 ;
        RECT 80.100 52.800 81.000 53.100 ;
        RECT 75.300 51.800 76.200 52.200 ;
        RECT 78.700 51.800 79.400 52.200 ;
        RECT 75.300 51.100 75.700 51.800 ;
        RECT 78.700 51.100 79.100 51.800 ;
        RECT 80.100 51.100 80.500 52.800 ;
        RECT 82.200 52.400 82.600 53.200 ;
        RECT 83.100 52.200 83.400 53.800 ;
        RECT 85.000 53.600 85.400 53.800 ;
        RECT 84.700 53.100 86.500 53.300 ;
        RECT 87.100 53.200 87.400 53.800 ;
        RECT 83.000 51.100 83.400 52.200 ;
        RECT 84.600 53.000 86.600 53.100 ;
        RECT 84.600 51.100 85.000 53.000 ;
        RECT 86.200 51.400 86.600 53.000 ;
        RECT 87.000 51.700 87.400 53.200 ;
        RECT 87.800 51.400 88.200 53.100 ;
        RECT 88.600 52.800 89.000 53.200 ;
        RECT 89.500 53.100 89.800 54.900 ;
        RECT 91.000 54.800 91.400 54.900 ;
        RECT 92.600 54.800 93.400 55.200 ;
        RECT 90.200 53.800 90.600 54.600 ;
        RECT 94.200 54.200 94.500 55.800 ;
        RECT 93.700 54.100 94.500 54.200 ;
        RECT 93.600 53.900 94.500 54.100 ;
        RECT 95.100 54.200 95.400 55.800 ;
        RECT 97.400 55.400 97.800 56.200 ;
        RECT 98.200 55.900 100.200 56.200 ;
        RECT 100.600 55.900 101.000 59.900 ;
        RECT 104.300 57.200 104.700 59.900 ;
        RECT 106.200 57.900 106.600 59.900 ;
        RECT 106.300 57.800 106.600 57.900 ;
        RECT 107.800 57.900 108.200 59.900 ;
        RECT 107.800 57.800 108.100 57.900 ;
        RECT 106.300 57.500 108.100 57.800 ;
        RECT 103.800 56.800 104.700 57.200 ;
        RECT 105.000 56.800 105.400 57.200 ;
        RECT 104.300 56.200 104.700 56.800 ;
        RECT 105.100 56.200 105.400 56.800 ;
        RECT 106.300 56.200 106.600 57.500 ;
        RECT 107.000 56.400 107.400 57.200 ;
        RECT 109.400 56.200 109.800 59.900 ;
        RECT 111.000 56.200 111.400 59.900 ;
        RECT 104.300 55.900 104.800 56.200 ;
        RECT 105.100 55.900 105.800 56.200 ;
        RECT 98.600 55.200 99.000 55.400 ;
        RECT 100.600 55.200 100.900 55.900 ;
        RECT 96.200 54.800 97.000 55.200 ;
        RECT 98.200 54.900 99.000 55.200 ;
        RECT 99.800 54.900 101.000 55.200 ;
        RECT 98.200 54.800 98.600 54.900 ;
        RECT 95.100 54.100 95.900 54.200 ;
        RECT 95.100 53.900 96.000 54.100 ;
        RECT 88.700 52.400 89.100 52.800 ;
        RECT 86.200 51.100 88.200 51.400 ;
        RECT 89.400 51.100 89.800 53.100 ;
        RECT 93.600 51.100 94.000 53.900 ;
        RECT 95.600 52.100 96.000 53.900 ;
        RECT 99.000 53.800 99.400 54.600 ;
        RECT 99.800 53.100 100.100 54.900 ;
        RECT 100.600 54.800 101.000 54.900 ;
        RECT 101.400 55.100 101.800 55.200 ;
        RECT 103.800 55.100 104.200 55.200 ;
        RECT 101.400 54.800 104.200 55.100 ;
        RECT 103.800 54.400 104.200 54.800 ;
        RECT 104.500 54.200 104.800 55.900 ;
        RECT 105.400 55.800 105.800 55.900 ;
        RECT 106.200 55.800 106.600 56.200 ;
        RECT 106.300 54.200 106.600 55.800 ;
        RECT 108.600 55.400 109.000 56.200 ;
        RECT 109.400 55.900 111.400 56.200 ;
        RECT 111.800 55.900 112.200 59.900 ;
        RECT 113.400 57.900 113.800 59.900 ;
        RECT 113.500 57.800 113.800 57.900 ;
        RECT 115.000 57.900 115.400 59.900 ;
        RECT 115.800 57.900 116.200 59.900 ;
        RECT 115.000 57.800 115.300 57.900 ;
        RECT 113.500 57.500 115.300 57.800 ;
        RECT 114.200 56.400 114.600 57.200 ;
        RECT 115.000 56.200 115.300 57.500 ;
        RECT 115.900 57.800 116.200 57.900 ;
        RECT 117.400 57.900 117.800 59.900 ;
        RECT 117.400 57.800 117.700 57.900 ;
        RECT 115.900 57.500 117.700 57.800 ;
        RECT 115.900 56.200 116.200 57.500 ;
        RECT 116.600 56.400 117.000 57.200 ;
        RECT 119.000 56.200 119.400 59.900 ;
        RECT 120.600 56.200 121.000 59.900 ;
        RECT 109.800 55.200 110.200 55.400 ;
        RECT 111.800 55.200 112.100 55.900 ;
        RECT 112.600 55.400 113.000 56.200 ;
        RECT 115.000 55.800 115.400 56.200 ;
        RECT 115.800 55.800 116.200 56.200 ;
        RECT 107.400 54.800 108.200 55.200 ;
        RECT 109.400 54.900 110.200 55.200 ;
        RECT 111.000 54.900 112.200 55.200 ;
        RECT 109.400 54.800 109.800 54.900 ;
        RECT 103.000 54.100 103.400 54.200 ;
        RECT 103.000 53.800 103.800 54.100 ;
        RECT 104.500 53.800 105.800 54.200 ;
        RECT 106.300 54.100 107.100 54.200 ;
        RECT 106.300 53.900 107.200 54.100 ;
        RECT 103.400 53.600 103.800 53.800 ;
        RECT 96.600 52.100 97.000 52.200 ;
        RECT 95.600 51.800 97.000 52.100 ;
        RECT 95.600 51.100 96.000 51.800 ;
        RECT 99.800 51.100 100.200 53.100 ;
        RECT 100.600 52.800 101.000 53.200 ;
        RECT 103.100 53.100 104.900 53.300 ;
        RECT 105.400 53.100 105.700 53.800 ;
        RECT 106.800 53.100 107.200 53.900 ;
        RECT 107.800 53.800 108.200 54.200 ;
        RECT 110.200 53.800 110.600 54.600 ;
        RECT 107.800 53.100 108.100 53.800 ;
        RECT 103.000 53.000 105.000 53.100 ;
        RECT 100.500 52.400 100.900 52.800 ;
        RECT 103.000 51.100 103.400 53.000 ;
        RECT 104.600 51.100 105.000 53.000 ;
        RECT 105.400 51.100 105.800 53.100 ;
        RECT 106.800 52.800 108.100 53.100 ;
        RECT 111.000 53.100 111.300 54.900 ;
        RECT 111.800 54.800 112.200 54.900 ;
        RECT 113.400 54.800 114.200 55.200 ;
        RECT 115.000 54.200 115.300 55.800 ;
        RECT 114.500 54.100 115.300 54.200 ;
        RECT 114.400 53.900 115.300 54.100 ;
        RECT 115.900 54.200 116.200 55.800 ;
        RECT 118.200 55.400 118.600 56.200 ;
        RECT 119.000 55.900 121.000 56.200 ;
        RECT 121.400 55.900 121.800 59.900 ;
        RECT 122.200 57.900 122.600 59.900 ;
        RECT 122.300 57.800 122.600 57.900 ;
        RECT 123.800 57.900 124.200 59.900 ;
        RECT 123.800 57.800 124.100 57.900 ;
        RECT 122.300 57.500 124.100 57.800 ;
        RECT 122.300 56.200 122.600 57.500 ;
        RECT 123.800 57.200 124.100 57.500 ;
        RECT 123.000 56.400 123.400 57.200 ;
        RECT 123.800 56.800 124.200 57.200 ;
        RECT 119.400 55.200 119.800 55.400 ;
        RECT 121.400 55.200 121.700 55.900 ;
        RECT 122.200 55.800 122.600 56.200 ;
        RECT 117.000 54.800 117.800 55.200 ;
        RECT 119.000 54.900 119.800 55.200 ;
        RECT 120.600 54.900 121.800 55.200 ;
        RECT 119.000 54.800 119.400 54.900 ;
        RECT 115.900 54.100 116.700 54.200 ;
        RECT 115.900 53.900 117.700 54.100 ;
        RECT 106.800 51.100 107.200 52.800 ;
        RECT 111.000 51.100 111.400 53.100 ;
        RECT 111.800 52.800 112.200 53.200 ;
        RECT 111.700 52.400 112.100 52.800 ;
        RECT 114.400 52.200 114.800 53.900 ;
        RECT 116.400 53.800 117.700 53.900 ;
        RECT 119.800 53.800 120.200 54.600 ;
        RECT 114.400 51.800 115.400 52.200 ;
        RECT 114.400 51.100 114.800 51.800 ;
        RECT 116.400 51.100 116.800 53.800 ;
        RECT 117.400 53.200 117.700 53.800 ;
        RECT 117.400 52.800 117.800 53.200 ;
        RECT 120.600 53.100 120.900 54.900 ;
        RECT 121.400 54.800 121.800 54.900 ;
        RECT 122.300 54.200 122.600 55.800 ;
        RECT 124.600 55.400 125.000 56.200 ;
        RECT 125.400 55.900 125.800 59.900 ;
        RECT 126.200 56.200 126.600 59.900 ;
        RECT 127.800 56.200 128.200 59.900 ;
        RECT 129.900 58.200 130.300 59.900 ;
        RECT 129.400 57.800 130.300 58.200 ;
        RECT 131.800 57.900 132.200 59.900 ;
        RECT 126.200 55.900 128.200 56.200 ;
        RECT 129.900 56.200 130.300 57.800 ;
        RECT 131.900 57.800 132.200 57.900 ;
        RECT 133.400 57.900 133.800 59.900 ;
        RECT 135.800 57.900 136.200 59.900 ;
        RECT 133.400 57.800 133.700 57.900 ;
        RECT 131.900 57.500 133.700 57.800 ;
        RECT 135.900 57.800 136.200 57.900 ;
        RECT 137.400 57.900 137.800 59.900 ;
        RECT 137.400 57.800 137.700 57.900 ;
        RECT 135.900 57.500 137.700 57.800 ;
        RECT 130.600 56.800 131.000 57.200 ;
        RECT 130.700 56.200 131.000 56.800 ;
        RECT 131.900 56.200 132.200 57.500 ;
        RECT 132.600 57.100 133.000 57.200 ;
        RECT 136.600 57.100 137.000 57.200 ;
        RECT 132.600 56.800 137.000 57.100 ;
        RECT 132.600 56.400 133.000 56.800 ;
        RECT 136.600 56.400 137.000 56.800 ;
        RECT 137.400 56.200 137.700 57.500 ;
        RECT 129.900 55.900 130.400 56.200 ;
        RECT 130.700 55.900 131.400 56.200 ;
        RECT 125.500 55.200 125.800 55.900 ;
        RECT 127.400 55.200 127.800 55.400 ;
        RECT 123.400 54.800 124.200 55.200 ;
        RECT 125.400 54.900 126.600 55.200 ;
        RECT 127.400 54.900 128.200 55.200 ;
        RECT 125.400 54.800 125.800 54.900 ;
        RECT 122.300 54.100 123.100 54.200 ;
        RECT 122.300 53.900 123.200 54.100 ;
        RECT 120.600 51.100 121.000 53.100 ;
        RECT 121.400 52.800 121.800 53.200 ;
        RECT 121.300 52.400 121.700 52.800 ;
        RECT 122.800 51.100 123.200 53.900 ;
        RECT 126.300 53.200 126.600 54.900 ;
        RECT 127.800 54.800 128.200 54.900 ;
        RECT 127.000 53.800 127.400 54.600 ;
        RECT 129.400 54.400 129.800 55.200 ;
        RECT 130.100 54.200 130.400 55.900 ;
        RECT 131.000 55.800 131.400 55.900 ;
        RECT 131.800 55.800 132.200 56.200 ;
        RECT 131.900 54.200 132.200 55.800 ;
        RECT 134.200 56.100 134.600 56.200 ;
        RECT 135.000 56.100 135.400 56.200 ;
        RECT 134.200 55.800 135.400 56.100 ;
        RECT 134.200 55.400 134.600 55.800 ;
        RECT 135.000 55.400 135.400 55.800 ;
        RECT 137.400 55.800 137.800 56.200 ;
        RECT 133.000 54.800 133.800 55.200 ;
        RECT 135.800 54.800 136.600 55.200 ;
        RECT 137.400 54.200 137.700 55.800 ;
        RECT 128.600 54.100 129.000 54.200 ;
        RECT 128.600 53.800 129.400 54.100 ;
        RECT 130.100 53.800 131.400 54.200 ;
        RECT 131.900 54.100 132.700 54.200 ;
        RECT 136.900 54.100 137.700 54.200 ;
        RECT 131.900 53.900 132.800 54.100 ;
        RECT 129.000 53.600 129.400 53.800 ;
        RECT 125.400 52.800 125.800 53.200 ;
        RECT 125.500 52.400 125.900 52.800 ;
        RECT 126.200 51.100 126.600 53.200 ;
        RECT 128.700 53.100 130.500 53.300 ;
        RECT 131.000 53.100 131.300 53.800 ;
        RECT 128.600 53.000 130.600 53.100 ;
        RECT 128.600 51.100 129.000 53.000 ;
        RECT 130.200 51.100 130.600 53.000 ;
        RECT 131.000 51.100 131.400 53.100 ;
        RECT 132.400 52.200 132.800 53.900 ;
        RECT 131.800 51.800 132.800 52.200 ;
        RECT 132.400 51.100 132.800 51.800 ;
        RECT 136.800 53.900 137.700 54.100 ;
        RECT 136.800 52.200 137.200 53.900 ;
        RECT 138.200 53.400 138.600 54.200 ;
        RECT 139.000 54.100 139.400 59.900 ;
        RECT 139.800 55.800 140.200 56.600 ;
        RECT 139.800 54.800 140.200 55.200 ;
        RECT 139.800 54.100 140.100 54.800 ;
        RECT 139.000 53.800 140.100 54.100 ;
        RECT 139.000 53.100 139.400 53.800 ;
        RECT 139.000 52.800 139.900 53.100 ;
        RECT 136.800 51.800 137.800 52.200 ;
        RECT 136.800 51.100 137.200 51.800 ;
        RECT 139.500 51.100 139.900 52.800 ;
        RECT 140.600 51.100 141.000 59.900 ;
        RECT 142.200 56.200 142.600 59.900 ;
        RECT 143.000 56.200 143.400 56.300 ;
        RECT 144.400 56.200 145.200 59.900 ;
        RECT 142.200 55.900 143.400 56.200 ;
        RECT 144.200 55.900 145.200 56.200 ;
        RECT 146.300 56.200 146.700 56.300 ;
        RECT 147.000 56.200 147.400 59.900 ;
        RECT 149.100 57.200 149.500 59.900 ;
        RECT 148.600 56.800 149.500 57.200 ;
        RECT 149.800 56.800 150.200 57.200 ;
        RECT 146.300 55.900 147.400 56.200 ;
        RECT 149.100 56.200 149.500 56.800 ;
        RECT 149.900 56.200 150.200 56.800 ;
        RECT 149.100 55.900 149.600 56.200 ;
        RECT 149.900 55.900 150.600 56.200 ;
        RECT 144.200 55.200 144.500 55.900 ;
        RECT 146.300 55.600 146.600 55.900 ;
        RECT 144.900 55.300 146.600 55.600 ;
        RECT 144.900 55.200 145.300 55.300 ;
        RECT 143.800 54.900 144.500 55.200 ;
        RECT 146.000 54.900 146.400 55.000 ;
        RECT 143.800 54.800 144.700 54.900 ;
        RECT 144.200 54.600 144.700 54.800 ;
        RECT 141.400 54.100 141.800 54.200 ;
        RECT 142.200 54.100 143.000 54.200 ;
        RECT 141.400 53.800 143.000 54.100 ;
        RECT 143.600 53.800 144.000 54.200 ;
        RECT 141.400 53.400 141.800 53.800 ;
        RECT 143.700 53.600 144.000 53.800 ;
        RECT 143.000 53.400 143.400 53.500 ;
        RECT 142.200 53.100 143.400 53.400 ;
        RECT 143.700 53.200 144.100 53.600 ;
        RECT 142.200 51.100 142.600 53.100 ;
        RECT 144.400 52.900 144.700 54.600 ;
        RECT 145.100 54.600 146.400 54.900 ;
        RECT 145.100 54.300 145.400 54.600 ;
        RECT 148.600 54.400 149.000 55.200 ;
        RECT 145.000 53.900 145.400 54.300 ;
        RECT 149.300 54.200 149.600 55.900 ;
        RECT 150.200 55.800 150.600 55.900 ;
        RECT 146.600 54.100 147.400 54.200 ;
        RECT 145.700 53.800 147.400 54.100 ;
        RECT 147.800 54.100 148.200 54.200 ;
        RECT 147.800 53.800 148.600 54.100 ;
        RECT 149.300 53.800 150.600 54.200 ;
        RECT 145.700 53.600 146.000 53.800 ;
        RECT 148.200 53.600 148.600 53.800 ;
        RECT 145.000 53.300 146.000 53.600 ;
        RECT 146.300 53.400 146.700 53.500 ;
        RECT 145.000 53.200 145.800 53.300 ;
        RECT 146.300 53.100 147.400 53.400 ;
        RECT 147.900 53.100 149.700 53.300 ;
        RECT 150.200 53.100 150.500 53.800 ;
        RECT 144.400 52.200 145.200 52.900 ;
        RECT 144.400 51.800 145.800 52.200 ;
        RECT 144.400 51.100 145.200 51.800 ;
        RECT 147.000 51.100 147.400 53.100 ;
        RECT 147.800 53.000 149.800 53.100 ;
        RECT 147.800 51.100 148.200 53.000 ;
        RECT 149.400 51.100 149.800 53.000 ;
        RECT 150.200 51.100 150.600 53.100 ;
        RECT 1.900 48.200 2.300 49.900 ;
        RECT 1.400 47.900 2.300 48.200 ;
        RECT 3.000 47.900 3.400 49.900 ;
        RECT 5.200 48.100 6.000 49.900 ;
        RECT 1.400 46.100 1.800 47.900 ;
        RECT 3.000 47.600 4.200 47.900 ;
        RECT 3.800 47.500 4.200 47.600 ;
        RECT 5.200 46.400 5.500 48.100 ;
        RECT 7.800 47.900 8.200 49.900 ;
        RECT 8.600 47.900 9.000 49.900 ;
        RECT 9.400 48.000 9.800 49.900 ;
        RECT 11.000 48.000 11.400 49.900 ;
        RECT 9.400 47.900 11.400 48.000 ;
        RECT 11.800 47.900 12.200 49.900 ;
        RECT 14.000 48.100 14.800 49.900 ;
        RECT 7.100 47.600 8.200 47.900 ;
        RECT 7.100 47.500 7.500 47.600 ;
        RECT 8.700 47.200 9.000 47.900 ;
        RECT 9.500 47.700 11.300 47.900 ;
        RECT 11.800 47.600 13.000 47.900 ;
        RECT 12.600 47.500 13.000 47.600 ;
        RECT 13.300 47.400 13.700 47.800 ;
        RECT 10.600 47.200 11.000 47.400 ;
        RECT 13.300 47.200 13.600 47.400 ;
        RECT 5.800 46.700 6.200 47.100 ;
        RECT 8.600 46.800 9.900 47.200 ;
        RECT 10.600 46.900 11.400 47.200 ;
        RECT 11.000 46.800 11.400 46.900 ;
        RECT 11.800 46.800 12.600 47.200 ;
        RECT 13.200 46.800 13.600 47.200 ;
        RECT 14.000 47.100 14.300 48.100 ;
        RECT 16.600 47.900 17.000 49.900 ;
        RECT 14.600 47.400 15.400 47.800 ;
        RECT 15.700 47.600 17.000 47.900 ;
        RECT 15.700 47.500 16.100 47.600 ;
        RECT 17.400 47.500 17.800 49.900 ;
        RECT 19.600 49.200 20.000 49.900 ;
        RECT 19.000 48.900 20.000 49.200 ;
        RECT 21.800 48.900 22.200 49.900 ;
        RECT 23.900 49.200 24.500 49.900 ;
        RECT 23.800 48.900 24.500 49.200 ;
        RECT 19.000 48.500 19.400 48.900 ;
        RECT 21.800 48.600 22.100 48.900 ;
        RECT 19.800 48.200 20.200 48.600 ;
        RECT 20.700 48.300 22.100 48.600 ;
        RECT 23.800 48.500 24.200 48.900 ;
        RECT 20.700 48.200 21.100 48.300 ;
        RECT 16.200 47.100 17.000 47.200 ;
        RECT 14.000 46.800 14.500 47.100 ;
        RECT 15.900 47.000 17.000 47.100 ;
        RECT 5.000 46.200 5.500 46.400 ;
        RECT 3.000 46.100 3.400 46.200 ;
        RECT 1.400 45.800 3.400 46.100 ;
        RECT 4.600 46.100 5.500 46.200 ;
        RECT 5.900 46.400 6.200 46.700 ;
        RECT 5.900 46.100 7.200 46.400 ;
        RECT 4.600 45.800 5.300 46.100 ;
        RECT 6.800 46.000 7.200 46.100 ;
        RECT 1.400 41.100 1.800 45.800 ;
        RECT 5.000 45.100 5.300 45.800 ;
        RECT 5.700 45.700 6.100 45.800 ;
        RECT 5.700 45.400 7.400 45.700 ;
        RECT 7.100 45.100 7.400 45.400 ;
        RECT 8.600 45.100 9.000 45.200 ;
        RECT 9.600 45.100 9.900 46.800 ;
        RECT 10.200 46.100 10.600 46.600 ;
        RECT 11.800 46.100 12.100 46.800 ;
        RECT 14.200 46.200 14.500 46.800 ;
        RECT 14.800 46.800 17.000 47.000 ;
        RECT 17.800 47.100 18.600 47.200 ;
        RECT 19.900 47.100 20.200 48.200 ;
        RECT 24.700 47.700 25.100 47.800 ;
        RECT 26.200 47.700 26.600 49.900 ;
        RECT 24.700 47.400 26.600 47.700 ;
        RECT 27.800 47.600 28.200 49.900 ;
        RECT 29.400 47.600 29.800 49.900 ;
        RECT 31.000 47.600 31.400 49.900 ;
        RECT 32.600 47.600 33.000 49.900 ;
        RECT 35.000 48.900 35.400 49.900 ;
        RECT 34.200 48.100 34.600 48.200 ;
        RECT 35.000 48.100 35.300 48.900 ;
        RECT 34.200 47.800 35.300 48.100 ;
        RECT 22.700 47.100 23.100 47.200 ;
        RECT 17.800 46.800 23.300 47.100 ;
        RECT 14.800 46.700 16.200 46.800 ;
        RECT 19.300 46.700 19.700 46.800 ;
        RECT 14.800 46.600 15.200 46.700 ;
        RECT 18.500 46.200 18.900 46.300 ;
        RECT 19.800 46.200 20.200 46.300 ;
        RECT 23.000 46.200 23.300 46.800 ;
        RECT 23.800 46.400 24.200 46.500 ;
        RECT 10.200 45.800 12.100 46.100 ;
        RECT 13.400 46.100 13.800 46.200 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 15.500 46.100 15.900 46.200 ;
        RECT 13.400 45.800 14.600 46.100 ;
        RECT 15.100 45.800 15.900 46.100 ;
        RECT 18.500 45.900 21.000 46.200 ;
        RECT 20.600 45.800 21.000 45.900 ;
        RECT 23.000 45.800 23.400 46.200 ;
        RECT 23.800 46.100 25.700 46.400 ;
        RECT 25.300 46.000 25.700 46.100 ;
        RECT 14.200 45.100 14.500 45.800 ;
        RECT 15.100 45.700 15.500 45.800 ;
        RECT 17.400 45.500 20.200 45.600 ;
        RECT 17.400 45.400 20.300 45.500 ;
        RECT 17.400 45.300 22.300 45.400 ;
        RECT 3.000 44.800 4.200 45.100 ;
        RECT 5.000 44.800 6.000 45.100 ;
        RECT 3.000 41.100 3.400 44.800 ;
        RECT 3.800 44.700 4.200 44.800 ;
        RECT 5.200 44.200 6.000 44.800 ;
        RECT 7.100 44.800 8.200 45.100 ;
        RECT 8.600 44.800 9.300 45.100 ;
        RECT 9.600 44.800 10.100 45.100 ;
        RECT 7.100 44.700 7.500 44.800 ;
        RECT 5.200 43.800 6.600 44.200 ;
        RECT 5.200 41.100 6.000 43.800 ;
        RECT 7.800 41.100 8.200 44.800 ;
        RECT 9.000 44.200 9.300 44.800 ;
        RECT 9.000 43.800 9.400 44.200 ;
        RECT 9.700 41.100 10.100 44.800 ;
        RECT 11.800 44.800 13.000 45.100 ;
        RECT 11.800 41.100 12.200 44.800 ;
        RECT 12.600 44.700 13.000 44.800 ;
        RECT 14.000 41.100 14.800 45.100 ;
        RECT 15.700 44.800 17.000 45.100 ;
        RECT 15.700 44.700 16.100 44.800 ;
        RECT 16.600 41.100 17.000 44.800 ;
        RECT 17.400 41.100 17.800 45.300 ;
        RECT 19.900 45.100 22.300 45.300 ;
        RECT 19.000 44.500 21.700 44.800 ;
        RECT 19.000 44.400 19.400 44.500 ;
        RECT 21.300 44.400 21.700 44.500 ;
        RECT 22.000 44.500 22.300 45.100 ;
        RECT 23.000 45.200 23.300 45.800 ;
        RECT 24.500 45.700 24.900 45.800 ;
        RECT 26.200 45.700 26.600 47.400 ;
        RECT 24.500 45.400 26.600 45.700 ;
        RECT 27.000 47.200 28.200 47.600 ;
        RECT 28.700 47.200 29.800 47.600 ;
        RECT 30.300 47.200 31.400 47.600 ;
        RECT 32.100 47.200 33.000 47.600 ;
        RECT 35.000 47.200 35.300 47.800 ;
        RECT 35.800 47.800 36.200 48.600 ;
        RECT 36.600 47.900 37.000 49.900 ;
        RECT 38.700 48.400 39.100 49.900 ;
        RECT 38.700 47.900 39.400 48.400 ;
        RECT 39.800 48.000 40.200 49.900 ;
        RECT 41.400 48.000 41.800 49.900 ;
        RECT 39.800 47.900 41.800 48.000 ;
        RECT 42.200 47.900 42.600 49.900 ;
        RECT 36.700 47.800 37.000 47.900 ;
        RECT 27.000 45.800 27.400 47.200 ;
        RECT 28.700 46.900 29.100 47.200 ;
        RECT 30.300 46.900 30.700 47.200 ;
        RECT 32.100 46.900 32.500 47.200 ;
        RECT 27.800 46.500 29.100 46.900 ;
        RECT 29.500 46.500 30.700 46.900 ;
        RECT 31.200 46.500 32.500 46.900 ;
        RECT 28.700 45.800 29.100 46.500 ;
        RECT 30.300 45.800 30.700 46.500 ;
        RECT 32.100 45.800 32.500 46.500 ;
        RECT 35.000 46.800 35.400 47.200 ;
        RECT 35.800 47.100 36.100 47.800 ;
        RECT 36.700 47.600 37.600 47.800 ;
        RECT 36.700 47.500 38.800 47.600 ;
        RECT 37.300 47.300 38.800 47.500 ;
        RECT 38.400 47.200 38.800 47.300 ;
        RECT 36.600 47.100 37.000 47.200 ;
        RECT 35.800 46.800 37.000 47.100 ;
        RECT 37.600 46.900 38.000 47.000 ;
        RECT 27.000 45.400 28.200 45.800 ;
        RECT 28.700 45.400 29.800 45.800 ;
        RECT 30.300 45.400 31.400 45.800 ;
        RECT 32.100 45.400 33.000 45.800 ;
        RECT 34.200 45.400 34.600 46.200 ;
        RECT 23.000 44.900 24.200 45.200 ;
        RECT 22.700 44.500 23.100 44.600 ;
        RECT 22.000 44.200 23.100 44.500 ;
        RECT 23.900 44.400 24.200 44.900 ;
        RECT 23.900 44.000 24.600 44.400 ;
        RECT 20.700 43.700 21.100 43.800 ;
        RECT 22.100 43.700 22.500 43.800 ;
        RECT 19.000 43.100 19.400 43.500 ;
        RECT 20.700 43.400 22.500 43.700 ;
        RECT 21.800 43.100 22.100 43.400 ;
        RECT 23.800 43.100 24.200 43.500 ;
        RECT 19.000 42.800 20.000 43.100 ;
        RECT 19.600 41.100 20.000 42.800 ;
        RECT 21.800 41.100 22.200 43.100 ;
        RECT 23.900 41.100 24.500 43.100 ;
        RECT 26.200 41.100 26.600 45.400 ;
        RECT 27.800 41.100 28.200 45.400 ;
        RECT 29.400 41.100 29.800 45.400 ;
        RECT 31.000 41.100 31.400 45.400 ;
        RECT 32.600 41.100 33.000 45.400 ;
        RECT 35.000 45.100 35.300 46.800 ;
        RECT 36.600 46.400 37.000 46.800 ;
        RECT 37.500 46.600 38.000 46.900 ;
        RECT 37.500 46.200 37.800 46.600 ;
        RECT 37.400 45.800 37.800 46.200 ;
        RECT 38.400 45.500 38.700 47.200 ;
        RECT 39.100 46.200 39.400 47.900 ;
        RECT 39.900 47.700 41.700 47.900 ;
        RECT 40.200 47.200 40.600 47.400 ;
        RECT 42.200 47.200 42.500 47.900 ;
        RECT 39.800 46.900 40.600 47.200 ;
        RECT 39.800 46.800 40.200 46.900 ;
        RECT 41.300 46.800 42.600 47.200 ;
        RECT 39.000 46.100 39.400 46.200 ;
        RECT 39.800 46.100 40.200 46.200 ;
        RECT 39.000 45.800 40.200 46.100 ;
        RECT 40.600 45.800 41.000 46.600 ;
        RECT 37.500 45.200 38.700 45.500 ;
        RECT 34.500 44.700 35.400 45.100 ;
        RECT 34.500 41.100 34.900 44.700 ;
        RECT 37.500 43.100 37.800 45.200 ;
        RECT 39.100 45.100 39.400 45.800 ;
        RECT 41.300 45.100 41.600 46.800 ;
        RECT 42.200 46.200 42.500 46.800 ;
        RECT 42.200 45.800 42.600 46.200 ;
        RECT 42.200 45.100 42.600 45.200 ;
        RECT 37.400 41.100 37.800 43.100 ;
        RECT 39.000 41.100 39.400 45.100 ;
        RECT 41.100 44.800 41.600 45.100 ;
        RECT 41.900 44.800 42.600 45.100 ;
        RECT 41.100 41.100 41.500 44.800 ;
        RECT 41.900 44.200 42.200 44.800 ;
        RECT 41.800 43.800 42.200 44.200 ;
        RECT 43.000 41.100 43.400 49.900 ;
        RECT 45.400 48.900 45.800 49.900 ;
        RECT 43.800 47.800 44.200 48.600 ;
        RECT 44.600 47.800 45.000 48.600 ;
        RECT 43.800 47.100 44.100 47.800 ;
        RECT 45.500 47.200 45.800 48.900 ;
        RECT 47.100 48.200 47.500 48.600 ;
        RECT 46.200 48.100 46.600 48.200 ;
        RECT 47.000 48.100 47.400 48.200 ;
        RECT 46.200 47.800 47.400 48.100 ;
        RECT 47.800 47.900 48.200 49.900 ;
        RECT 44.600 47.100 45.000 47.200 ;
        RECT 43.800 46.800 45.000 47.100 ;
        RECT 45.400 47.100 45.800 47.200 ;
        RECT 47.000 47.100 47.400 47.200 ;
        RECT 45.400 46.800 47.400 47.100 ;
        RECT 45.500 45.100 45.800 46.800 ;
        RECT 46.200 45.400 46.600 46.200 ;
        RECT 47.000 46.100 47.400 46.200 ;
        RECT 47.900 46.100 48.200 47.900 ;
        RECT 51.800 47.900 52.200 49.900 ;
        RECT 54.000 49.200 54.800 49.900 ;
        RECT 53.400 48.800 54.800 49.200 ;
        RECT 54.000 48.100 54.800 48.800 ;
        RECT 51.800 47.600 53.000 47.900 ;
        RECT 52.600 47.500 53.000 47.600 ;
        RECT 53.300 47.400 53.700 47.800 ;
        RECT 53.300 47.200 53.600 47.400 ;
        RECT 48.600 46.400 49.000 47.200 ;
        RECT 51.800 47.100 52.600 47.200 ;
        RECT 49.400 46.800 52.600 47.100 ;
        RECT 53.200 46.800 53.600 47.200 ;
        RECT 54.000 47.100 54.300 48.100 ;
        RECT 56.600 47.900 57.000 49.900 ;
        RECT 54.600 47.400 55.400 47.800 ;
        RECT 55.700 47.600 57.000 47.900 ;
        RECT 55.700 47.500 56.100 47.600 ;
        RECT 57.400 47.500 57.800 49.900 ;
        RECT 59.600 49.200 60.000 49.900 ;
        RECT 59.000 48.900 60.000 49.200 ;
        RECT 61.800 48.900 62.200 49.900 ;
        RECT 63.900 49.200 64.500 49.900 ;
        RECT 63.800 48.900 64.500 49.200 ;
        RECT 59.000 48.500 59.400 48.900 ;
        RECT 61.800 48.600 62.100 48.900 ;
        RECT 59.800 48.200 60.200 48.600 ;
        RECT 60.700 48.300 62.100 48.600 ;
        RECT 63.800 48.500 64.200 48.900 ;
        RECT 60.700 48.200 61.100 48.300 ;
        RECT 56.200 47.100 57.000 47.200 ;
        RECT 54.000 46.800 54.500 47.100 ;
        RECT 55.900 47.000 57.000 47.100 ;
        RECT 49.400 46.200 49.700 46.800 ;
        RECT 54.200 46.200 54.500 46.800 ;
        RECT 54.800 46.800 57.000 47.000 ;
        RECT 57.800 47.100 58.600 47.200 ;
        RECT 59.900 47.100 60.200 48.200 ;
        RECT 64.700 47.700 65.100 47.800 ;
        RECT 66.200 47.700 66.600 49.900 ;
        RECT 64.700 47.400 66.600 47.700 ;
        RECT 67.800 47.600 68.200 49.900 ;
        RECT 69.400 47.600 69.800 49.900 ;
        RECT 71.000 47.600 71.400 49.900 ;
        RECT 72.600 47.600 73.000 49.900 ;
        RECT 75.000 48.900 75.400 49.900 ;
        RECT 74.200 47.800 74.600 48.600 ;
        RECT 62.700 47.100 63.100 47.200 ;
        RECT 57.800 46.800 63.300 47.100 ;
        RECT 54.800 46.700 56.200 46.800 ;
        RECT 59.300 46.700 59.700 46.800 ;
        RECT 54.800 46.600 55.200 46.700 ;
        RECT 58.500 46.200 58.900 46.300 ;
        RECT 59.800 46.200 60.200 46.300 ;
        RECT 63.000 46.200 63.300 46.800 ;
        RECT 63.800 46.400 64.200 46.500 ;
        RECT 49.400 46.100 49.800 46.200 ;
        RECT 47.000 45.800 48.200 46.100 ;
        RECT 49.000 45.800 49.800 46.100 ;
        RECT 54.200 45.800 54.600 46.200 ;
        RECT 55.500 46.100 55.900 46.200 ;
        RECT 55.100 45.800 55.900 46.100 ;
        RECT 58.500 45.900 61.000 46.200 ;
        RECT 60.600 45.800 61.000 45.900 ;
        RECT 63.000 45.800 63.400 46.200 ;
        RECT 63.800 46.100 65.700 46.400 ;
        RECT 65.300 46.000 65.700 46.100 ;
        RECT 47.100 45.100 47.400 45.800 ;
        RECT 49.000 45.600 49.400 45.800 ;
        RECT 54.200 45.100 54.500 45.800 ;
        RECT 55.100 45.700 55.500 45.800 ;
        RECT 57.400 45.500 60.200 45.600 ;
        RECT 57.400 45.400 60.300 45.500 ;
        RECT 57.400 45.300 62.300 45.400 ;
        RECT 45.400 44.700 46.300 45.100 ;
        RECT 45.900 41.100 46.300 44.700 ;
        RECT 47.000 41.100 47.400 45.100 ;
        RECT 47.800 44.800 49.800 45.100 ;
        RECT 47.800 41.100 48.200 44.800 ;
        RECT 49.400 41.100 49.800 44.800 ;
        RECT 51.800 44.800 53.000 45.100 ;
        RECT 51.800 41.100 52.200 44.800 ;
        RECT 52.600 44.700 53.000 44.800 ;
        RECT 54.000 41.100 54.800 45.100 ;
        RECT 55.700 44.800 57.000 45.100 ;
        RECT 55.700 44.700 56.100 44.800 ;
        RECT 56.600 41.100 57.000 44.800 ;
        RECT 57.400 41.100 57.800 45.300 ;
        RECT 59.900 45.100 62.300 45.300 ;
        RECT 59.000 44.500 61.700 44.800 ;
        RECT 59.000 44.400 59.400 44.500 ;
        RECT 61.300 44.400 61.700 44.500 ;
        RECT 62.000 44.500 62.300 45.100 ;
        RECT 63.000 45.200 63.300 45.800 ;
        RECT 64.500 45.700 64.900 45.800 ;
        RECT 66.200 45.700 66.600 47.400 ;
        RECT 64.500 45.400 66.600 45.700 ;
        RECT 67.000 47.200 68.200 47.600 ;
        RECT 68.700 47.200 69.800 47.600 ;
        RECT 70.300 47.200 71.400 47.600 ;
        RECT 72.100 47.200 73.000 47.600 ;
        RECT 75.100 47.200 75.400 48.900 ;
        RECT 76.600 47.900 77.000 49.900 ;
        RECT 77.400 48.000 77.800 49.900 ;
        RECT 79.000 48.000 79.400 49.900 ;
        RECT 77.400 47.900 79.400 48.000 ;
        RECT 76.700 47.200 77.000 47.900 ;
        RECT 77.500 47.700 79.300 47.900 ;
        RECT 78.600 47.200 79.000 47.400 ;
        RECT 67.000 45.800 67.400 47.200 ;
        RECT 68.700 46.900 69.100 47.200 ;
        RECT 70.300 46.900 70.700 47.200 ;
        RECT 72.100 46.900 72.500 47.200 ;
        RECT 67.800 46.500 69.100 46.900 ;
        RECT 69.500 46.500 70.700 46.900 ;
        RECT 71.200 46.500 72.500 46.900 ;
        RECT 75.000 46.800 75.400 47.200 ;
        RECT 76.600 46.800 77.900 47.200 ;
        RECT 78.600 47.100 79.400 47.200 ;
        RECT 79.800 47.100 80.200 49.900 ;
        RECT 80.600 47.800 81.000 48.600 ;
        RECT 81.400 47.900 81.800 49.900 ;
        RECT 82.200 48.000 82.600 49.900 ;
        RECT 83.800 48.000 84.200 49.900 ;
        RECT 82.200 47.900 84.200 48.000 ;
        RECT 81.500 47.200 81.800 47.900 ;
        RECT 82.300 47.700 84.100 47.900 ;
        RECT 83.400 47.200 83.800 47.400 ;
        RECT 78.600 46.900 80.200 47.100 ;
        RECT 79.000 46.800 80.200 46.900 ;
        RECT 81.400 46.800 82.700 47.200 ;
        RECT 83.400 46.900 84.200 47.200 ;
        RECT 83.800 46.800 84.200 46.900 ;
        RECT 84.600 46.800 85.000 47.600 ;
        RECT 85.400 47.100 85.800 49.900 ;
        RECT 87.000 48.800 87.400 49.900 ;
        RECT 89.400 48.900 89.800 49.900 ;
        RECT 86.200 47.800 86.600 48.600 ;
        RECT 87.100 47.200 87.400 48.800 ;
        RECT 88.600 48.100 89.000 48.600 ;
        RECT 87.800 47.800 89.000 48.100 ;
        RECT 89.500 47.200 89.800 48.900 ;
        RECT 91.000 47.600 91.400 49.900 ;
        RECT 92.600 48.200 93.000 49.900 ;
        RECT 92.600 47.900 93.100 48.200 ;
        RECT 91.000 47.300 92.300 47.600 ;
        RECT 85.400 46.800 86.500 47.100 ;
        RECT 87.000 46.800 87.400 47.200 ;
        RECT 89.400 46.800 89.800 47.200 ;
        RECT 68.700 45.800 69.100 46.500 ;
        RECT 70.300 45.800 70.700 46.500 ;
        RECT 72.100 45.800 72.500 46.500 ;
        RECT 67.000 45.400 68.200 45.800 ;
        RECT 68.700 45.400 69.800 45.800 ;
        RECT 70.300 45.400 71.400 45.800 ;
        RECT 72.100 45.400 73.000 45.800 ;
        RECT 63.000 44.900 64.200 45.200 ;
        RECT 62.700 44.500 63.100 44.600 ;
        RECT 62.000 44.200 63.100 44.500 ;
        RECT 63.900 44.400 64.200 44.900 ;
        RECT 63.900 44.000 64.600 44.400 ;
        RECT 60.700 43.700 61.100 43.800 ;
        RECT 62.100 43.700 62.500 43.800 ;
        RECT 59.000 43.100 59.400 43.500 ;
        RECT 60.700 43.400 62.500 43.700 ;
        RECT 61.800 43.100 62.100 43.400 ;
        RECT 63.800 43.100 64.200 43.500 ;
        RECT 59.000 42.800 60.000 43.100 ;
        RECT 59.600 41.100 60.000 42.800 ;
        RECT 61.800 41.100 62.200 43.100 ;
        RECT 63.900 41.100 64.500 43.100 ;
        RECT 66.200 41.100 66.600 45.400 ;
        RECT 67.800 41.100 68.200 45.400 ;
        RECT 69.400 41.100 69.800 45.400 ;
        RECT 71.000 41.100 71.400 45.400 ;
        RECT 72.600 41.100 73.000 45.400 ;
        RECT 75.100 45.100 75.400 46.800 ;
        RECT 75.800 46.100 76.200 46.200 ;
        RECT 75.800 45.800 76.900 46.100 ;
        RECT 75.800 45.400 76.200 45.800 ;
        RECT 76.600 45.200 76.900 45.800 ;
        RECT 77.600 45.200 77.900 46.800 ;
        RECT 78.200 45.800 78.600 46.600 ;
        RECT 76.600 45.100 77.000 45.200 ;
        RECT 75.000 44.700 75.900 45.100 ;
        RECT 76.600 44.800 77.300 45.100 ;
        RECT 77.600 44.800 78.600 45.200 ;
        RECT 75.500 44.200 75.900 44.700 ;
        RECT 77.000 44.200 77.300 44.800 ;
        RECT 75.500 43.800 76.200 44.200 ;
        RECT 77.000 43.800 77.400 44.200 ;
        RECT 75.500 41.100 75.900 43.800 ;
        RECT 77.700 41.100 78.100 44.800 ;
        RECT 79.800 41.100 80.200 46.800 ;
        RECT 81.400 45.100 81.800 45.200 ;
        RECT 82.400 45.100 82.700 46.800 ;
        RECT 83.000 45.800 83.400 46.600 ;
        RECT 81.400 44.800 82.100 45.100 ;
        RECT 82.400 44.800 82.900 45.100 ;
        RECT 81.800 44.200 82.100 44.800 ;
        RECT 81.800 43.800 82.200 44.200 ;
        RECT 82.500 41.100 82.900 44.800 ;
        RECT 85.400 41.100 85.800 46.800 ;
        RECT 86.200 46.200 86.500 46.800 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 87.100 45.100 87.400 46.800 ;
        RECT 87.800 45.400 88.200 46.200 ;
        RECT 88.600 46.100 89.000 46.200 ;
        RECT 89.500 46.100 89.800 46.800 ;
        RECT 91.100 46.200 91.500 46.600 ;
        RECT 88.600 45.800 89.800 46.100 ;
        RECT 89.500 45.100 89.800 45.800 ;
        RECT 90.200 45.400 90.600 46.200 ;
        RECT 91.000 45.800 91.500 46.200 ;
        RECT 92.000 46.500 92.300 47.300 ;
        RECT 92.800 47.200 93.100 47.900 ;
        RECT 92.600 46.800 93.100 47.200 ;
        RECT 94.200 46.800 94.600 47.600 ;
        RECT 92.000 46.100 92.500 46.500 ;
        RECT 92.000 45.100 92.300 46.100 ;
        RECT 92.800 45.100 93.100 46.800 ;
        RECT 87.000 44.700 87.900 45.100 ;
        RECT 89.400 44.700 90.300 45.100 ;
        RECT 87.500 41.100 87.900 44.700 ;
        RECT 89.900 41.100 90.300 44.700 ;
        RECT 91.000 44.800 92.300 45.100 ;
        RECT 91.000 41.100 91.400 44.800 ;
        RECT 92.600 44.600 93.100 45.100 ;
        RECT 95.000 45.100 95.400 49.900 ;
        RECT 95.800 47.900 96.200 49.900 ;
        RECT 96.600 48.000 97.000 49.900 ;
        RECT 98.200 48.000 98.600 49.900 ;
        RECT 96.600 47.900 98.600 48.000 ;
        RECT 99.800 48.900 100.200 49.900 ;
        RECT 95.900 47.200 96.200 47.900 ;
        RECT 96.700 47.700 98.500 47.900 ;
        RECT 97.800 47.200 98.200 47.400 ;
        RECT 99.800 47.200 100.100 48.900 ;
        RECT 100.600 47.800 101.000 48.600 ;
        RECT 103.100 48.200 103.500 48.600 ;
        RECT 103.000 47.800 103.400 48.200 ;
        RECT 103.800 47.900 104.200 49.900 ;
        RECT 95.800 46.800 97.100 47.200 ;
        RECT 97.800 46.900 98.600 47.200 ;
        RECT 96.800 46.200 97.100 46.800 ;
        RECT 98.200 46.800 98.600 46.900 ;
        RECT 99.800 46.800 100.200 47.200 ;
        RECT 95.800 45.800 96.200 46.200 ;
        RECT 96.600 45.800 97.100 46.200 ;
        RECT 97.400 45.800 97.800 46.600 ;
        RECT 98.200 46.100 98.500 46.800 ;
        RECT 99.000 46.100 99.400 46.200 ;
        RECT 98.200 45.800 99.400 46.100 ;
        RECT 95.800 45.200 96.100 45.800 ;
        RECT 95.800 45.100 96.200 45.200 ;
        RECT 96.800 45.100 97.100 45.800 ;
        RECT 99.000 45.400 99.400 45.800 ;
        RECT 99.800 45.100 100.100 46.800 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 103.900 46.100 104.200 47.900 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 106.200 47.100 106.600 49.900 ;
        RECT 107.000 47.800 107.400 48.600 ;
        RECT 107.800 48.000 108.200 49.900 ;
        RECT 109.400 48.000 109.800 49.900 ;
        RECT 107.800 47.900 109.800 48.000 ;
        RECT 110.200 47.900 110.600 49.900 ;
        RECT 111.000 48.000 111.400 49.900 ;
        RECT 112.600 48.000 113.000 49.900 ;
        RECT 111.000 47.900 113.000 48.000 ;
        RECT 113.400 47.900 113.800 49.900 ;
        RECT 107.900 47.700 109.700 47.900 ;
        RECT 108.200 47.200 108.600 47.400 ;
        RECT 110.200 47.200 110.500 47.900 ;
        RECT 111.100 47.700 112.900 47.900 ;
        RECT 111.400 47.200 111.800 47.400 ;
        RECT 113.400 47.200 113.700 47.900 ;
        RECT 114.200 47.800 114.600 48.600 ;
        RECT 104.600 46.800 106.600 47.100 ;
        RECT 107.800 46.900 108.600 47.200 ;
        RECT 107.800 46.800 108.200 46.900 ;
        RECT 109.300 46.800 110.600 47.200 ;
        RECT 111.000 46.900 111.800 47.200 ;
        RECT 111.000 46.800 111.400 46.900 ;
        RECT 112.500 46.800 113.800 47.200 ;
        RECT 104.600 46.400 105.000 46.800 ;
        RECT 105.400 46.100 105.800 46.200 ;
        RECT 103.000 45.800 104.200 46.100 ;
        RECT 105.000 45.800 105.800 46.100 ;
        RECT 103.100 45.100 103.400 45.800 ;
        RECT 105.000 45.600 105.400 45.800 ;
        RECT 95.000 44.800 96.500 45.100 ;
        RECT 96.800 44.800 97.300 45.100 ;
        RECT 92.600 41.100 93.000 44.600 ;
        RECT 95.000 41.100 95.400 44.800 ;
        RECT 96.200 44.200 96.500 44.800 ;
        RECT 96.200 43.800 96.600 44.200 ;
        RECT 96.900 41.100 97.300 44.800 ;
        RECT 99.300 44.700 100.200 45.100 ;
        RECT 99.300 42.200 99.700 44.700 ;
        RECT 99.300 41.800 100.200 42.200 ;
        RECT 99.300 41.100 99.700 41.800 ;
        RECT 103.000 41.100 103.400 45.100 ;
        RECT 103.800 44.800 105.800 45.100 ;
        RECT 103.800 41.100 104.200 44.800 ;
        RECT 105.400 41.100 105.800 44.800 ;
        RECT 106.200 41.100 106.600 46.800 ;
        RECT 107.000 46.100 107.400 46.200 ;
        RECT 108.600 46.100 109.000 46.600 ;
        RECT 107.000 45.800 109.000 46.100 ;
        RECT 109.300 45.100 109.600 46.800 ;
        RECT 111.800 45.800 112.200 46.600 ;
        RECT 112.500 46.200 112.800 46.800 ;
        RECT 112.500 45.800 113.000 46.200 ;
        RECT 110.200 45.100 110.600 45.200 ;
        RECT 112.500 45.100 112.800 45.800 ;
        RECT 113.400 45.100 113.800 45.200 ;
        RECT 114.200 45.100 114.600 45.200 ;
        RECT 109.100 44.800 109.600 45.100 ;
        RECT 109.900 44.800 110.600 45.100 ;
        RECT 112.300 44.800 112.800 45.100 ;
        RECT 113.100 44.800 114.600 45.100 ;
        RECT 109.100 42.200 109.500 44.800 ;
        RECT 109.900 44.200 110.200 44.800 ;
        RECT 109.800 43.800 110.200 44.200 ;
        RECT 108.600 41.800 109.500 42.200 ;
        RECT 109.100 41.100 109.500 41.800 ;
        RECT 112.300 41.100 112.700 44.800 ;
        RECT 113.100 44.200 113.400 44.800 ;
        RECT 113.000 43.800 113.400 44.200 ;
        RECT 115.000 41.100 115.400 49.900 ;
        RECT 115.900 48.200 116.300 48.600 ;
        RECT 115.800 47.800 116.200 48.200 ;
        RECT 116.600 47.900 117.000 49.900 ;
        RECT 115.800 46.100 116.200 46.200 ;
        RECT 116.700 46.100 117.000 47.900 ;
        RECT 117.400 46.400 117.800 47.200 ;
        RECT 120.800 47.100 121.200 49.900 ;
        RECT 120.800 46.900 121.700 47.100 ;
        RECT 120.900 46.800 121.700 46.900 ;
        RECT 122.200 46.800 122.600 47.600 ;
        RECT 118.200 46.100 118.600 46.200 ;
        RECT 115.800 45.800 117.000 46.100 ;
        RECT 117.800 45.800 118.600 46.100 ;
        RECT 119.800 45.800 120.600 46.200 ;
        RECT 115.900 45.100 116.200 45.800 ;
        RECT 117.800 45.600 118.200 45.800 ;
        RECT 115.800 41.100 116.200 45.100 ;
        RECT 116.600 44.800 118.600 45.100 ;
        RECT 119.000 44.800 119.400 45.600 ;
        RECT 121.400 45.200 121.700 46.800 ;
        RECT 121.400 44.800 121.800 45.200 ;
        RECT 116.600 41.100 117.000 44.800 ;
        RECT 118.200 41.100 118.600 44.800 ;
        RECT 120.600 43.800 121.000 44.600 ;
        RECT 121.400 43.500 121.700 44.800 ;
        RECT 119.900 43.200 121.700 43.500 ;
        RECT 119.900 43.100 120.200 43.200 ;
        RECT 119.800 41.100 120.200 43.100 ;
        RECT 121.400 43.100 121.700 43.200 ;
        RECT 121.400 41.100 121.800 43.100 ;
        RECT 123.000 41.100 123.400 49.900 ;
        RECT 125.400 47.900 125.800 49.900 ;
        RECT 126.100 48.200 126.500 48.600 ;
        RECT 124.600 46.400 125.000 47.200 ;
        RECT 123.800 46.100 124.200 46.200 ;
        RECT 125.400 46.100 125.700 47.900 ;
        RECT 126.200 47.800 126.600 48.200 ;
        RECT 127.000 48.000 127.400 49.900 ;
        RECT 128.600 48.000 129.000 49.900 ;
        RECT 127.000 47.900 129.000 48.000 ;
        RECT 129.400 47.900 129.800 49.900 ;
        RECT 127.100 47.700 128.900 47.900 ;
        RECT 127.400 47.200 127.800 47.400 ;
        RECT 129.400 47.200 129.700 47.900 ;
        RECT 127.000 46.900 127.800 47.200 ;
        RECT 127.000 46.800 127.400 46.900 ;
        RECT 128.500 46.800 129.800 47.200 ;
        RECT 130.800 47.100 131.200 49.900 ;
        RECT 133.500 48.200 133.900 48.600 ;
        RECT 133.400 47.800 133.800 48.200 ;
        RECT 134.200 47.900 134.600 49.900 ;
        RECT 137.400 48.900 137.800 49.900 ;
        RECT 130.300 46.900 131.200 47.100 ;
        RECT 130.300 46.800 131.100 46.900 ;
        RECT 126.200 46.100 126.600 46.200 ;
        RECT 123.800 45.800 124.600 46.100 ;
        RECT 125.400 45.800 126.600 46.100 ;
        RECT 127.800 45.800 128.200 46.600 ;
        RECT 128.500 46.200 128.800 46.800 ;
        RECT 128.500 45.800 129.000 46.200 ;
        RECT 124.200 45.600 124.600 45.800 ;
        RECT 126.200 45.100 126.500 45.800 ;
        RECT 128.500 45.100 128.800 45.800 ;
        RECT 130.300 45.200 130.600 46.800 ;
        RECT 131.400 45.800 132.200 46.200 ;
        RECT 133.400 46.100 133.800 46.200 ;
        RECT 134.300 46.100 134.600 47.900 ;
        RECT 136.600 47.800 137.000 48.600 ;
        RECT 137.500 47.800 137.800 48.900 ;
        RECT 139.000 47.900 139.400 49.900 ;
        RECT 141.100 48.200 141.500 49.900 ;
        RECT 137.500 47.500 138.700 47.800 ;
        RECT 135.000 46.400 135.400 47.200 ;
        RECT 137.400 46.800 137.900 47.200 ;
        RECT 137.600 46.400 138.000 46.800 ;
        RECT 135.800 46.100 136.200 46.200 ;
        RECT 133.400 45.800 134.600 46.100 ;
        RECT 135.400 45.800 136.200 46.100 ;
        RECT 138.400 46.000 138.700 47.500 ;
        RECT 139.100 46.200 139.400 47.900 ;
        RECT 140.600 47.900 141.500 48.200 ;
        RECT 139.800 46.800 140.200 47.600 ;
        RECT 129.400 45.100 129.800 45.200 ;
        RECT 123.800 44.800 125.800 45.100 ;
        RECT 123.800 41.100 124.200 44.800 ;
        RECT 125.400 41.100 125.800 44.800 ;
        RECT 126.200 41.100 126.600 45.100 ;
        RECT 128.300 44.800 128.800 45.100 ;
        RECT 129.100 44.800 129.800 45.100 ;
        RECT 130.200 44.800 130.600 45.200 ;
        RECT 132.600 44.800 133.000 45.600 ;
        RECT 133.500 45.100 133.800 45.800 ;
        RECT 135.400 45.600 135.800 45.800 ;
        RECT 138.300 45.700 138.700 46.000 ;
        RECT 139.000 45.800 139.400 46.200 ;
        RECT 136.600 45.600 138.700 45.700 ;
        RECT 136.600 45.400 138.600 45.600 ;
        RECT 128.300 41.100 128.700 44.800 ;
        RECT 129.100 44.200 129.400 44.800 ;
        RECT 129.000 43.800 129.400 44.200 ;
        RECT 130.300 43.500 130.600 44.800 ;
        RECT 131.000 43.800 131.400 44.600 ;
        RECT 130.300 43.200 132.100 43.500 ;
        RECT 130.300 43.100 130.600 43.200 ;
        RECT 130.200 41.100 130.600 43.100 ;
        RECT 131.800 43.100 132.100 43.200 ;
        RECT 131.800 41.100 132.200 43.100 ;
        RECT 133.400 41.100 133.800 45.100 ;
        RECT 134.200 44.800 136.200 45.100 ;
        RECT 134.200 41.100 134.600 44.800 ;
        RECT 135.800 41.100 136.200 44.800 ;
        RECT 136.600 41.100 137.000 45.400 ;
        RECT 139.100 45.100 139.400 45.800 ;
        RECT 139.800 45.800 140.200 46.200 ;
        RECT 140.600 46.100 141.000 47.900 ;
        RECT 144.000 47.100 144.400 49.900 ;
        RECT 146.200 48.900 146.600 49.900 ;
        RECT 145.400 47.800 145.800 48.600 ;
        RECT 146.300 47.200 146.600 48.900 ;
        RECT 147.800 47.900 148.200 49.900 ;
        RECT 149.900 48.400 150.300 49.900 ;
        RECT 149.900 47.900 150.600 48.400 ;
        RECT 147.900 47.800 148.200 47.900 ;
        RECT 147.900 47.600 148.800 47.800 ;
        RECT 147.900 47.500 150.000 47.600 ;
        RECT 148.500 47.300 150.000 47.500 ;
        RECT 149.600 47.200 150.000 47.300 ;
        RECT 144.000 46.900 144.900 47.100 ;
        RECT 144.100 46.800 144.900 46.900 ;
        RECT 146.200 46.800 146.600 47.200 ;
        RECT 147.000 47.100 147.400 47.200 ;
        RECT 147.800 47.100 148.200 47.200 ;
        RECT 147.000 46.800 148.200 47.100 ;
        RECT 148.800 46.900 149.200 47.000 ;
        RECT 140.600 45.800 142.600 46.100 ;
        RECT 143.000 45.800 143.800 46.200 ;
        RECT 139.800 45.100 140.100 45.800 ;
        RECT 138.700 44.800 140.100 45.100 ;
        RECT 138.700 41.100 139.100 44.800 ;
        RECT 140.600 41.100 141.000 45.800 ;
        RECT 141.400 44.400 141.800 45.200 ;
        RECT 142.200 44.800 142.600 45.800 ;
        RECT 144.600 45.200 144.900 46.800 ;
        RECT 144.600 44.800 145.000 45.200 ;
        RECT 146.300 45.100 146.600 46.800 ;
        RECT 147.000 46.100 147.400 46.200 ;
        RECT 147.800 46.100 148.200 46.800 ;
        RECT 148.700 46.600 149.200 46.900 ;
        RECT 148.700 46.200 149.000 46.600 ;
        RECT 147.000 45.800 148.200 46.100 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 147.000 45.400 147.400 45.800 ;
        RECT 149.600 45.500 149.900 47.200 ;
        RECT 150.300 46.200 150.600 47.900 ;
        RECT 150.200 45.800 150.600 46.200 ;
        RECT 148.700 45.200 149.900 45.500 ;
        RECT 143.800 43.800 144.200 44.600 ;
        RECT 144.600 43.500 144.900 44.800 ;
        RECT 146.200 44.700 147.100 45.100 ;
        RECT 143.100 43.200 144.900 43.500 ;
        RECT 143.100 43.100 143.400 43.200 ;
        RECT 143.000 41.100 143.400 43.100 ;
        RECT 144.600 43.100 144.900 43.200 ;
        RECT 146.700 44.100 147.100 44.700 ;
        RECT 147.800 44.100 148.200 44.200 ;
        RECT 146.700 43.800 148.200 44.100 ;
        RECT 144.600 41.100 145.000 43.100 ;
        RECT 146.700 41.100 147.100 43.800 ;
        RECT 148.700 43.100 149.000 45.200 ;
        RECT 150.300 45.100 150.600 45.800 ;
        RECT 148.600 41.100 149.000 43.100 ;
        RECT 150.200 41.100 150.600 45.100 ;
        RECT 0.600 36.200 1.000 39.900 ;
        RECT 1.500 36.200 1.900 36.300 ;
        RECT 0.600 35.900 1.900 36.200 ;
        RECT 2.800 35.900 3.600 39.900 ;
        RECT 4.600 36.200 5.000 36.300 ;
        RECT 5.400 36.200 5.800 39.900 ;
        RECT 4.600 35.900 5.800 36.200 ;
        RECT 2.100 35.200 2.500 35.300 ;
        RECT 3.100 35.200 3.400 35.900 ;
        RECT 1.700 34.900 2.500 35.200 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 1.700 34.800 2.100 34.900 ;
        RECT 3.000 34.800 4.200 35.100 ;
        RECT 3.100 34.200 3.400 34.800 ;
        RECT 3.100 33.900 3.600 34.200 ;
        RECT 1.500 33.400 1.900 33.500 ;
        RECT 0.600 33.100 1.900 33.400 ;
        RECT 2.200 33.200 3.000 33.600 ;
        RECT 0.600 31.100 1.000 33.100 ;
        RECT 3.300 32.900 3.600 33.900 ;
        RECT 4.000 33.800 4.400 34.200 ;
        RECT 4.000 33.600 4.300 33.800 ;
        RECT 3.900 33.200 4.300 33.600 ;
        RECT 4.600 33.400 5.000 33.500 ;
        RECT 4.600 33.100 5.800 33.400 ;
        RECT 2.800 31.100 3.600 32.900 ;
        RECT 5.400 31.100 5.800 33.100 ;
        RECT 7.000 33.100 7.400 39.900 ;
        RECT 7.800 36.100 8.200 36.600 ;
        RECT 8.600 36.100 9.000 39.900 ;
        RECT 10.600 36.800 11.000 37.200 ;
        RECT 10.600 36.200 10.900 36.800 ;
        RECT 11.300 36.200 11.700 39.900 ;
        RECT 7.800 35.800 9.000 36.100 ;
        RECT 10.200 35.900 10.900 36.200 ;
        RECT 11.200 35.900 11.700 36.200 ;
        RECT 13.400 36.200 13.800 39.900 ;
        RECT 14.200 36.200 14.600 36.300 ;
        RECT 13.400 35.900 14.600 36.200 ;
        RECT 15.600 36.200 16.400 39.900 ;
        RECT 17.300 36.200 17.700 36.300 ;
        RECT 18.200 36.200 18.600 39.900 ;
        RECT 15.600 35.900 17.000 36.200 ;
        RECT 17.300 35.900 18.600 36.200 ;
        RECT 10.200 35.800 10.600 35.900 ;
        RECT 7.000 32.800 7.900 33.100 ;
        RECT 7.500 31.100 7.900 32.800 ;
        RECT 8.600 31.100 9.000 35.800 ;
        RECT 11.200 34.200 11.500 35.900 ;
        RECT 15.800 35.800 17.000 35.900 ;
        RECT 15.800 35.200 16.100 35.800 ;
        RECT 19.000 35.700 19.400 39.900 ;
        RECT 21.200 38.200 21.600 39.900 ;
        RECT 20.600 37.900 21.600 38.200 ;
        RECT 23.400 37.900 23.800 39.900 ;
        RECT 25.500 37.900 26.100 39.900 ;
        RECT 20.600 37.500 21.000 37.900 ;
        RECT 23.400 37.600 23.700 37.900 ;
        RECT 22.300 37.300 24.100 37.600 ;
        RECT 25.400 37.500 25.800 37.900 ;
        RECT 22.300 37.200 22.700 37.300 ;
        RECT 23.700 37.200 24.100 37.300 ;
        RECT 20.600 36.500 21.000 36.600 ;
        RECT 22.900 36.500 23.300 36.600 ;
        RECT 20.600 36.200 23.300 36.500 ;
        RECT 23.600 36.500 24.700 36.800 ;
        RECT 23.600 35.900 23.900 36.500 ;
        RECT 24.300 36.400 24.700 36.500 ;
        RECT 25.500 36.600 26.200 37.000 ;
        RECT 25.500 36.100 25.800 36.600 ;
        RECT 21.500 35.700 23.900 35.900 ;
        RECT 19.000 35.600 23.900 35.700 ;
        RECT 24.600 35.800 25.800 36.100 ;
        RECT 19.000 35.500 21.900 35.600 ;
        RECT 19.000 35.400 21.800 35.500 ;
        RECT 16.700 35.200 17.100 35.300 ;
        RECT 11.800 35.100 12.200 35.200 ;
        RECT 11.800 34.800 13.700 35.100 ;
        RECT 11.800 34.400 12.200 34.800 ;
        RECT 13.400 34.200 13.700 34.800 ;
        RECT 15.800 34.800 16.200 35.200 ;
        RECT 16.700 34.900 17.500 35.200 ;
        RECT 22.200 35.100 22.600 35.200 ;
        RECT 17.100 34.800 17.500 34.900 ;
        RECT 20.100 34.800 22.600 35.100 ;
        RECT 15.800 34.200 16.100 34.800 ;
        RECT 20.100 34.700 20.500 34.800 ;
        RECT 21.400 34.700 21.800 34.800 ;
        RECT 10.200 33.800 11.500 34.200 ;
        RECT 12.600 34.100 13.000 34.200 ;
        RECT 12.200 33.800 13.000 34.100 ;
        RECT 13.400 33.800 14.200 34.200 ;
        RECT 14.800 33.800 15.200 34.200 ;
        RECT 10.300 33.100 10.600 33.800 ;
        RECT 12.200 33.600 12.600 33.800 ;
        RECT 14.900 33.600 15.200 33.800 ;
        RECT 15.600 33.900 16.100 34.200 ;
        RECT 16.400 34.300 16.800 34.400 ;
        RECT 16.400 34.200 17.800 34.300 ;
        RECT 20.900 34.200 21.300 34.300 ;
        RECT 24.600 34.200 24.900 35.800 ;
        RECT 27.800 35.600 28.200 39.900 ;
        RECT 26.100 35.300 28.200 35.600 ;
        RECT 28.600 35.700 29.000 39.900 ;
        RECT 30.800 38.200 31.200 39.900 ;
        RECT 30.200 37.900 31.200 38.200 ;
        RECT 33.000 37.900 33.400 39.900 ;
        RECT 35.100 37.900 35.700 39.900 ;
        RECT 30.200 37.500 30.600 37.900 ;
        RECT 33.000 37.600 33.300 37.900 ;
        RECT 31.900 37.300 33.700 37.600 ;
        RECT 35.000 37.500 35.400 37.900 ;
        RECT 31.900 37.200 32.300 37.300 ;
        RECT 33.300 37.200 33.700 37.300 ;
        RECT 30.200 36.500 30.600 36.600 ;
        RECT 32.500 36.500 32.900 36.600 ;
        RECT 30.200 36.200 32.900 36.500 ;
        RECT 33.200 36.500 34.300 36.800 ;
        RECT 33.200 35.900 33.500 36.500 ;
        RECT 33.900 36.400 34.300 36.500 ;
        RECT 35.100 36.600 35.800 37.000 ;
        RECT 35.100 36.100 35.400 36.600 ;
        RECT 31.100 35.700 33.500 35.900 ;
        RECT 28.600 35.600 33.500 35.700 ;
        RECT 34.200 35.800 35.400 36.100 ;
        RECT 28.600 35.500 31.500 35.600 ;
        RECT 28.600 35.400 31.400 35.500 ;
        RECT 26.100 35.200 26.500 35.300 ;
        RECT 26.900 34.900 27.300 35.000 ;
        RECT 25.400 34.600 27.300 34.900 ;
        RECT 25.400 34.500 25.800 34.600 ;
        RECT 16.400 34.000 18.600 34.200 ;
        RECT 17.500 33.900 18.600 34.000 ;
        RECT 14.200 33.400 14.600 33.500 ;
        RECT 11.100 33.100 12.900 33.300 ;
        RECT 13.400 33.100 14.600 33.400 ;
        RECT 14.900 33.200 15.300 33.600 ;
        RECT 10.200 31.100 10.600 33.100 ;
        RECT 11.000 33.000 13.000 33.100 ;
        RECT 11.000 31.100 11.400 33.000 ;
        RECT 12.600 31.100 13.000 33.000 ;
        RECT 13.400 31.100 13.800 33.100 ;
        RECT 15.600 32.900 15.900 33.900 ;
        RECT 17.800 33.800 18.600 33.900 ;
        RECT 19.400 33.900 24.900 34.200 ;
        RECT 19.400 33.800 20.200 33.900 ;
        RECT 16.200 33.200 17.000 33.600 ;
        RECT 17.300 33.400 17.700 33.500 ;
        RECT 17.300 33.100 18.600 33.400 ;
        RECT 15.600 31.100 16.400 32.900 ;
        RECT 18.200 31.100 18.600 33.100 ;
        RECT 19.000 31.100 19.400 33.500 ;
        RECT 21.500 33.200 21.800 33.900 ;
        RECT 24.300 33.800 24.700 33.900 ;
        RECT 27.800 33.600 28.200 35.300 ;
        RECT 30.500 34.200 30.900 34.300 ;
        RECT 34.200 34.200 34.500 35.800 ;
        RECT 37.400 35.600 37.800 39.900 ;
        RECT 35.700 35.300 37.800 35.600 ;
        RECT 35.700 35.200 36.100 35.300 ;
        RECT 36.500 34.900 36.900 35.000 ;
        RECT 35.000 34.600 36.900 34.900 ;
        RECT 35.000 34.500 35.400 34.600 ;
        RECT 29.000 33.900 34.500 34.200 ;
        RECT 29.000 33.800 29.800 33.900 ;
        RECT 26.300 33.300 28.200 33.600 ;
        RECT 26.300 33.200 26.700 33.300 ;
        RECT 20.600 32.100 21.000 32.500 ;
        RECT 21.400 32.400 21.800 33.200 ;
        RECT 22.300 32.700 22.700 32.800 ;
        RECT 22.300 32.400 23.700 32.700 ;
        RECT 23.400 32.100 23.700 32.400 ;
        RECT 25.400 32.100 25.800 32.500 ;
        RECT 20.600 31.800 21.600 32.100 ;
        RECT 21.200 31.100 21.600 31.800 ;
        RECT 23.400 31.100 23.800 32.100 ;
        RECT 25.400 31.800 26.100 32.100 ;
        RECT 25.500 31.100 26.100 31.800 ;
        RECT 27.800 31.100 28.200 33.300 ;
        RECT 28.600 31.100 29.000 33.500 ;
        RECT 31.100 33.200 31.400 33.900 ;
        RECT 33.900 33.800 34.300 33.900 ;
        RECT 37.400 33.600 37.800 35.300 ;
        RECT 35.900 33.300 37.800 33.600 ;
        RECT 35.900 33.200 36.300 33.300 ;
        RECT 30.200 32.100 30.600 32.500 ;
        RECT 31.000 32.400 31.400 33.200 ;
        RECT 31.900 32.700 32.300 32.800 ;
        RECT 31.900 32.400 33.300 32.700 ;
        RECT 33.000 32.100 33.300 32.400 ;
        RECT 35.000 32.100 35.400 32.500 ;
        RECT 30.200 31.800 31.200 32.100 ;
        RECT 30.800 31.100 31.200 31.800 ;
        RECT 33.000 31.100 33.400 32.100 ;
        RECT 35.000 31.800 35.700 32.100 ;
        RECT 35.100 31.100 35.700 31.800 ;
        RECT 37.400 31.100 37.800 33.300 ;
        RECT 38.200 31.100 38.600 39.900 ;
        RECT 39.800 36.200 40.200 39.900 ;
        RECT 40.600 36.200 41.000 36.300 ;
        RECT 39.800 35.900 41.000 36.200 ;
        RECT 42.000 36.200 42.800 39.900 ;
        RECT 43.700 36.200 44.100 36.300 ;
        RECT 44.600 36.200 45.000 39.900 ;
        RECT 42.000 35.900 43.400 36.200 ;
        RECT 43.700 35.900 45.000 36.200 ;
        RECT 42.200 35.800 43.400 35.900 ;
        RECT 45.400 35.800 45.800 36.600 ;
        RECT 42.200 35.200 42.500 35.800 ;
        RECT 43.100 35.200 43.500 35.300 ;
        RECT 42.200 34.800 42.600 35.200 ;
        RECT 43.100 34.900 43.900 35.200 ;
        RECT 43.500 34.800 43.900 34.900 ;
        RECT 42.200 34.200 42.500 34.800 ;
        RECT 39.800 34.100 40.600 34.200 ;
        RECT 39.000 33.800 40.600 34.100 ;
        RECT 41.200 33.800 41.600 34.200 ;
        RECT 39.000 33.200 39.300 33.800 ;
        RECT 41.300 33.600 41.600 33.800 ;
        RECT 42.000 33.900 42.500 34.200 ;
        RECT 42.800 34.300 43.200 34.400 ;
        RECT 42.800 34.200 44.200 34.300 ;
        RECT 42.800 34.000 45.000 34.200 ;
        RECT 43.900 33.900 45.000 34.000 ;
        RECT 40.600 33.400 41.000 33.500 ;
        RECT 39.000 32.400 39.400 33.200 ;
        RECT 39.800 33.100 41.000 33.400 ;
        RECT 41.300 33.200 41.700 33.600 ;
        RECT 39.800 31.100 40.200 33.100 ;
        RECT 42.000 32.900 42.300 33.900 ;
        RECT 44.200 33.800 45.000 33.900 ;
        RECT 42.600 33.200 43.400 33.600 ;
        RECT 43.700 33.400 44.100 33.500 ;
        RECT 43.700 33.100 45.000 33.400 ;
        RECT 46.200 33.100 46.600 39.900 ;
        RECT 49.400 36.200 49.800 39.900 ;
        RECT 51.600 39.200 52.400 39.900 ;
        RECT 51.600 38.800 53.000 39.200 ;
        RECT 50.300 36.200 50.700 36.300 ;
        RECT 49.400 35.900 50.700 36.200 ;
        RECT 51.600 35.900 52.400 38.800 ;
        RECT 53.400 36.200 53.800 36.300 ;
        RECT 54.200 36.200 54.600 39.900 ;
        RECT 53.400 35.900 54.600 36.200 ;
        RECT 50.900 35.200 51.300 35.300 ;
        RECT 51.900 35.200 52.200 35.900 ;
        RECT 55.000 35.700 55.400 39.900 ;
        RECT 57.200 38.200 57.600 39.900 ;
        RECT 56.600 37.900 57.600 38.200 ;
        RECT 59.400 37.900 59.800 39.900 ;
        RECT 61.500 37.900 62.100 39.900 ;
        RECT 56.600 37.500 57.000 37.900 ;
        RECT 59.400 37.600 59.700 37.900 ;
        RECT 58.300 37.300 60.100 37.600 ;
        RECT 61.400 37.500 61.800 37.900 ;
        RECT 58.300 37.200 58.700 37.300 ;
        RECT 59.700 37.200 60.100 37.300 ;
        RECT 56.600 36.500 57.000 36.600 ;
        RECT 58.900 36.500 59.300 36.600 ;
        RECT 56.600 36.200 59.300 36.500 ;
        RECT 59.600 36.500 60.700 36.800 ;
        RECT 59.600 35.900 59.900 36.500 ;
        RECT 60.300 36.400 60.700 36.500 ;
        RECT 61.500 36.600 62.200 37.000 ;
        RECT 61.500 36.100 61.800 36.600 ;
        RECT 57.500 35.700 59.900 35.900 ;
        RECT 55.000 35.600 59.900 35.700 ;
        RECT 60.600 35.800 61.800 36.100 ;
        RECT 55.000 35.500 57.900 35.600 ;
        RECT 55.000 35.400 57.800 35.500 ;
        RECT 50.500 34.900 51.300 35.200 ;
        RECT 50.500 34.800 50.900 34.900 ;
        RECT 51.800 34.800 52.200 35.200 ;
        RECT 58.200 35.100 58.600 35.200 ;
        RECT 51.200 34.300 51.600 34.400 ;
        RECT 50.200 34.200 51.600 34.300 ;
        RECT 47.000 33.400 47.400 34.200 ;
        RECT 48.600 34.100 49.000 34.200 ;
        RECT 49.400 34.100 51.600 34.200 ;
        RECT 48.600 34.000 51.600 34.100 ;
        RECT 51.900 34.200 52.200 34.800 ;
        RECT 56.100 34.800 58.600 35.100 ;
        RECT 56.100 34.700 56.500 34.800 ;
        RECT 56.900 34.200 57.300 34.300 ;
        RECT 60.600 34.200 60.900 35.800 ;
        RECT 63.800 35.600 64.200 39.900 ;
        RECT 62.100 35.300 64.200 35.600 ;
        RECT 64.600 35.700 65.000 39.900 ;
        RECT 66.800 38.200 67.200 39.900 ;
        RECT 66.200 37.900 67.200 38.200 ;
        RECT 69.000 37.900 69.400 39.900 ;
        RECT 71.100 37.900 71.700 39.900 ;
        RECT 66.200 37.500 66.600 37.900 ;
        RECT 69.000 37.600 69.300 37.900 ;
        RECT 67.900 37.300 69.700 37.600 ;
        RECT 71.000 37.500 71.400 37.900 ;
        RECT 67.900 37.200 68.300 37.300 ;
        RECT 69.300 37.200 69.700 37.300 ;
        RECT 66.200 36.500 66.600 36.600 ;
        RECT 68.500 36.500 68.900 36.600 ;
        RECT 66.200 36.200 68.900 36.500 ;
        RECT 69.200 36.500 70.300 36.800 ;
        RECT 69.200 35.900 69.500 36.500 ;
        RECT 69.900 36.400 70.300 36.500 ;
        RECT 71.100 36.600 71.800 37.000 ;
        RECT 71.100 36.100 71.400 36.600 ;
        RECT 67.100 35.700 69.500 35.900 ;
        RECT 64.600 35.600 69.500 35.700 ;
        RECT 70.200 35.800 71.400 36.100 ;
        RECT 64.600 35.500 67.500 35.600 ;
        RECT 64.600 35.400 67.400 35.500 ;
        RECT 62.100 35.200 62.500 35.300 ;
        RECT 62.900 34.900 63.300 35.000 ;
        RECT 61.400 34.600 63.300 34.900 ;
        RECT 61.400 34.500 61.800 34.600 ;
        RECT 48.600 33.900 50.500 34.000 ;
        RECT 51.900 33.900 52.400 34.200 ;
        RECT 48.600 33.800 50.200 33.900 ;
        RECT 50.300 33.400 50.700 33.500 ;
        RECT 42.000 31.100 42.800 32.900 ;
        RECT 44.600 31.100 45.000 33.100 ;
        RECT 45.700 32.800 46.600 33.100 ;
        RECT 49.400 33.100 50.700 33.400 ;
        RECT 51.000 33.200 51.800 33.600 ;
        RECT 45.700 31.100 46.100 32.800 ;
        RECT 49.400 31.100 49.800 33.100 ;
        RECT 52.100 32.900 52.400 33.900 ;
        RECT 52.800 33.800 53.200 34.200 ;
        RECT 53.800 33.800 54.600 34.200 ;
        RECT 55.400 33.900 60.900 34.200 ;
        RECT 55.400 33.800 56.200 33.900 ;
        RECT 52.800 33.600 53.100 33.800 ;
        RECT 52.700 33.200 53.100 33.600 ;
        RECT 53.400 33.400 53.800 33.500 ;
        RECT 53.400 33.100 54.600 33.400 ;
        RECT 51.600 31.100 52.400 32.900 ;
        RECT 54.200 31.100 54.600 33.100 ;
        RECT 55.000 31.100 55.400 33.500 ;
        RECT 57.500 33.200 57.800 33.900 ;
        RECT 60.300 33.800 60.900 33.900 ;
        RECT 56.600 32.100 57.000 32.500 ;
        RECT 57.400 32.400 57.800 33.200 ;
        RECT 60.600 33.200 60.900 33.800 ;
        RECT 63.800 33.600 64.200 35.300 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 65.700 34.800 68.200 35.100 ;
        RECT 65.700 34.700 66.100 34.800 ;
        RECT 67.000 34.700 67.400 34.800 ;
        RECT 66.500 34.200 66.900 34.300 ;
        RECT 70.200 34.200 70.500 35.800 ;
        RECT 73.400 35.600 73.800 39.900 ;
        RECT 71.700 35.300 73.800 35.600 ;
        RECT 71.700 35.200 72.100 35.300 ;
        RECT 72.500 34.900 72.900 35.000 ;
        RECT 71.000 34.600 72.900 34.900 ;
        RECT 71.000 34.500 71.400 34.600 ;
        RECT 65.000 33.900 70.500 34.200 ;
        RECT 65.000 33.800 65.800 33.900 ;
        RECT 62.300 33.300 64.200 33.600 ;
        RECT 62.300 33.200 62.700 33.300 ;
        RECT 60.600 32.800 61.000 33.200 ;
        RECT 58.300 32.700 58.700 32.800 ;
        RECT 58.300 32.400 59.700 32.700 ;
        RECT 59.400 32.100 59.700 32.400 ;
        RECT 61.400 32.100 61.800 32.500 ;
        RECT 56.600 31.800 57.600 32.100 ;
        RECT 57.200 31.100 57.600 31.800 ;
        RECT 59.400 31.100 59.800 32.100 ;
        RECT 61.400 31.800 62.100 32.100 ;
        RECT 61.500 31.100 62.100 31.800 ;
        RECT 63.800 31.100 64.200 33.300 ;
        RECT 64.600 31.100 65.000 33.500 ;
        RECT 67.100 32.800 67.400 33.900 ;
        RECT 69.900 33.800 70.300 33.900 ;
        RECT 73.400 33.600 73.800 35.300 ;
        RECT 75.000 35.100 75.400 39.900 ;
        RECT 76.900 36.300 77.300 39.900 ;
        RECT 76.900 35.900 77.800 36.300 ;
        RECT 76.600 35.100 77.000 35.600 ;
        RECT 75.000 34.800 77.000 35.100 ;
        RECT 71.900 33.300 73.800 33.600 ;
        RECT 74.200 33.400 74.600 34.200 ;
        RECT 71.900 33.200 72.300 33.300 ;
        RECT 66.200 32.100 66.600 32.500 ;
        RECT 67.000 32.400 67.400 32.800 ;
        RECT 67.900 32.700 68.300 32.800 ;
        RECT 67.900 32.400 69.300 32.700 ;
        RECT 69.000 32.100 69.300 32.400 ;
        RECT 71.000 32.100 71.400 32.500 ;
        RECT 66.200 31.800 67.200 32.100 ;
        RECT 66.800 31.100 67.200 31.800 ;
        RECT 69.000 31.100 69.400 32.100 ;
        RECT 71.000 31.800 71.700 32.100 ;
        RECT 71.100 31.100 71.700 31.800 ;
        RECT 73.400 31.100 73.800 33.300 ;
        RECT 75.000 31.100 75.400 34.800 ;
        RECT 77.400 34.200 77.700 35.900 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 76.600 33.100 77.000 33.200 ;
        RECT 77.400 33.100 77.700 33.800 ;
        RECT 76.600 32.800 77.700 33.100 ;
        RECT 77.400 32.100 77.700 32.800 ;
        RECT 78.200 32.400 78.600 33.200 ;
        RECT 79.000 32.400 79.400 33.200 ;
        RECT 77.400 31.100 77.800 32.100 ;
        RECT 79.800 31.100 80.200 39.900 ;
        RECT 81.900 36.200 82.300 39.900 ;
        RECT 82.600 36.800 83.000 37.200 ;
        RECT 82.700 36.200 83.000 36.800 ;
        RECT 84.100 36.300 84.500 39.900 ;
        RECT 86.600 36.800 87.000 37.200 ;
        RECT 81.900 35.900 82.400 36.200 ;
        RECT 82.700 35.900 83.400 36.200 ;
        RECT 84.100 35.900 85.000 36.300 ;
        RECT 86.600 36.200 86.900 36.800 ;
        RECT 87.300 36.200 87.700 39.900 ;
        RECT 89.800 36.800 90.200 37.200 ;
        RECT 89.800 36.200 90.100 36.800 ;
        RECT 90.500 36.200 90.900 39.900 ;
        RECT 86.200 35.900 86.900 36.200 ;
        RECT 87.200 35.900 87.700 36.200 ;
        RECT 89.400 35.900 90.100 36.200 ;
        RECT 90.400 35.900 90.900 36.200 ;
        RECT 81.400 34.400 81.800 35.200 ;
        RECT 82.100 34.200 82.400 35.900 ;
        RECT 83.000 35.800 83.400 35.900 ;
        RECT 83.800 34.800 84.200 35.600 ;
        RECT 84.600 34.200 84.900 35.900 ;
        RECT 86.200 35.800 86.600 35.900 ;
        RECT 87.200 34.200 87.500 35.900 ;
        RECT 89.400 35.800 89.800 35.900 ;
        RECT 87.800 34.400 88.200 35.200 ;
        RECT 90.400 34.200 90.700 35.900 ;
        RECT 91.000 34.400 91.400 35.200 ;
        RECT 91.800 34.800 92.200 35.200 ;
        RECT 80.600 34.100 81.000 34.200 ;
        RECT 80.600 33.800 81.400 34.100 ;
        RECT 82.100 33.800 83.400 34.200 ;
        RECT 84.600 33.800 85.000 34.200 ;
        RECT 86.200 33.800 87.500 34.200 ;
        RECT 88.600 34.100 89.000 34.200 ;
        RECT 88.200 33.800 89.000 34.100 ;
        RECT 89.400 33.800 90.700 34.200 ;
        RECT 91.800 34.200 92.100 34.800 ;
        RECT 91.800 34.100 92.200 34.200 ;
        RECT 92.600 34.100 93.000 39.900 ;
        RECT 94.200 36.200 94.600 39.900 ;
        RECT 95.800 36.400 96.200 39.900 ;
        RECT 94.200 35.900 95.500 36.200 ;
        RECT 95.800 35.900 96.300 36.400 ;
        RECT 98.700 36.200 99.100 39.900 ;
        RECT 99.400 36.800 99.800 37.200 ;
        RECT 99.500 36.200 99.800 36.800 ;
        RECT 93.400 35.100 93.800 35.200 ;
        RECT 94.200 35.100 94.700 35.200 ;
        RECT 93.400 34.800 94.700 35.100 ;
        RECT 94.300 34.400 94.700 34.800 ;
        RECT 95.200 34.900 95.500 35.900 ;
        RECT 95.200 34.500 95.700 34.900 ;
        RECT 91.400 33.800 93.000 34.100 ;
        RECT 81.000 33.600 81.400 33.800 ;
        RECT 80.700 33.100 82.500 33.300 ;
        RECT 83.000 33.100 83.300 33.800 ;
        RECT 80.600 33.000 82.600 33.100 ;
        RECT 80.600 31.100 81.000 33.000 ;
        RECT 82.200 31.100 82.600 33.000 ;
        RECT 83.000 31.100 83.400 33.100 ;
        RECT 84.600 32.200 84.900 33.800 ;
        RECT 85.400 32.400 85.800 33.200 ;
        RECT 86.300 33.100 86.600 33.800 ;
        RECT 88.200 33.600 88.600 33.800 ;
        RECT 87.100 33.100 88.900 33.300 ;
        RECT 89.500 33.200 89.800 33.800 ;
        RECT 91.400 33.600 91.800 33.800 ;
        RECT 84.600 31.100 85.000 32.200 ;
        RECT 86.200 31.100 86.600 33.100 ;
        RECT 87.000 33.000 89.000 33.100 ;
        RECT 87.000 31.100 87.400 33.000 ;
        RECT 88.600 31.100 89.000 33.000 ;
        RECT 89.400 31.100 89.800 33.200 ;
        RECT 90.300 33.100 92.100 33.300 ;
        RECT 90.200 33.000 92.200 33.100 ;
        RECT 90.200 31.100 90.600 33.000 ;
        RECT 91.800 31.100 92.200 33.000 ;
        RECT 92.600 31.100 93.000 33.800 ;
        RECT 95.200 33.700 95.500 34.500 ;
        RECT 96.000 34.200 96.300 35.900 ;
        RECT 98.200 35.800 99.200 36.200 ;
        RECT 99.500 36.100 100.200 36.200 ;
        RECT 102.200 36.100 102.600 36.600 ;
        RECT 99.500 35.900 102.600 36.100 ;
        RECT 99.800 35.800 102.600 35.900 ;
        RECT 97.400 35.100 97.800 35.200 ;
        RECT 98.200 35.100 98.600 35.200 ;
        RECT 97.400 34.800 98.600 35.100 ;
        RECT 98.200 34.400 98.600 34.800 ;
        RECT 98.900 34.200 99.200 35.800 ;
        RECT 95.800 33.800 96.300 34.200 ;
        RECT 97.400 34.100 97.800 34.200 ;
        RECT 97.400 33.800 98.200 34.100 ;
        RECT 98.900 33.800 100.200 34.200 ;
        RECT 102.200 34.100 102.600 34.200 ;
        RECT 103.000 34.100 103.400 39.900 ;
        RECT 104.600 35.100 105.000 35.200 ;
        RECT 105.400 35.100 105.800 39.900 ;
        RECT 106.200 35.900 106.600 39.900 ;
        RECT 107.000 36.200 107.400 39.900 ;
        RECT 108.600 36.200 109.000 39.900 ;
        RECT 110.200 37.900 110.600 39.900 ;
        RECT 110.300 37.800 110.600 37.900 ;
        RECT 111.800 37.900 112.200 39.900 ;
        RECT 111.800 37.800 112.100 37.900 ;
        RECT 110.300 37.500 112.100 37.800 ;
        RECT 111.000 36.400 111.400 37.200 ;
        RECT 111.800 36.200 112.100 37.500 ;
        RECT 113.900 36.200 114.300 39.900 ;
        RECT 114.600 36.800 115.000 37.200 ;
        RECT 114.700 36.200 115.000 36.800 ;
        RECT 107.000 35.900 109.000 36.200 ;
        RECT 106.300 35.200 106.600 35.900 ;
        RECT 109.400 35.400 109.800 36.200 ;
        RECT 111.800 35.800 112.200 36.200 ;
        RECT 113.900 35.900 114.400 36.200 ;
        RECT 114.700 35.900 115.400 36.200 ;
        RECT 115.800 35.900 116.200 39.900 ;
        RECT 116.600 36.200 117.000 39.900 ;
        RECT 118.200 36.200 118.600 39.900 ;
        RECT 116.600 35.900 118.600 36.200 ;
        RECT 108.200 35.200 108.600 35.400 ;
        RECT 104.600 34.800 105.800 35.100 ;
        RECT 106.200 34.900 107.400 35.200 ;
        RECT 108.200 34.900 109.000 35.200 ;
        RECT 106.200 34.800 106.600 34.900 ;
        RECT 102.200 33.800 103.400 34.100 ;
        RECT 94.200 33.400 95.500 33.700 ;
        RECT 93.400 32.400 93.800 33.200 ;
        RECT 94.200 31.100 94.600 33.400 ;
        RECT 96.000 33.100 96.300 33.800 ;
        RECT 97.800 33.600 98.200 33.800 ;
        RECT 97.500 33.100 99.300 33.300 ;
        RECT 99.800 33.100 100.100 33.800 ;
        RECT 103.000 33.100 103.400 33.800 ;
        RECT 103.800 33.400 104.200 34.200 ;
        RECT 95.800 32.800 96.300 33.100 ;
        RECT 97.400 33.000 99.400 33.100 ;
        RECT 95.800 31.100 96.200 32.800 ;
        RECT 97.400 31.100 97.800 33.000 ;
        RECT 99.000 31.100 99.400 33.000 ;
        RECT 99.800 31.100 100.200 33.100 ;
        RECT 102.500 32.800 103.400 33.100 ;
        RECT 102.500 31.100 102.900 32.800 ;
        RECT 104.600 32.400 105.000 33.200 ;
        RECT 105.400 33.100 105.800 34.800 ;
        RECT 107.100 33.200 107.400 34.900 ;
        RECT 108.600 34.800 109.000 34.900 ;
        RECT 110.200 34.800 111.000 35.200 ;
        RECT 111.800 35.100 112.100 35.800 ;
        RECT 112.600 35.100 113.000 35.200 ;
        RECT 111.800 34.800 113.000 35.100 ;
        RECT 107.800 33.800 108.200 34.600 ;
        RECT 111.800 34.200 112.100 34.800 ;
        RECT 113.400 34.400 113.800 35.200 ;
        RECT 114.100 34.200 114.400 35.900 ;
        RECT 115.000 35.800 115.400 35.900 ;
        RECT 115.900 35.200 116.200 35.900 ;
        RECT 119.000 35.800 119.400 36.600 ;
        RECT 117.800 35.200 118.200 35.400 ;
        RECT 115.800 34.900 117.000 35.200 ;
        RECT 117.800 35.100 118.600 35.200 ;
        RECT 119.000 35.100 119.400 35.200 ;
        RECT 117.800 34.900 119.400 35.100 ;
        RECT 115.800 34.800 116.200 34.900 ;
        RECT 111.300 34.100 112.100 34.200 ;
        RECT 111.200 33.900 112.100 34.100 ;
        RECT 112.600 34.100 113.000 34.200 ;
        RECT 106.200 33.100 106.600 33.200 ;
        RECT 105.400 32.800 106.600 33.100 ;
        RECT 105.400 31.100 105.800 32.800 ;
        RECT 106.300 32.400 106.700 32.800 ;
        RECT 107.000 31.100 107.400 33.200 ;
        RECT 111.200 31.100 111.600 33.900 ;
        RECT 112.600 33.800 113.400 34.100 ;
        RECT 114.100 33.800 115.400 34.200 ;
        RECT 113.000 33.600 113.400 33.800 ;
        RECT 112.700 33.100 114.500 33.300 ;
        RECT 115.000 33.100 115.300 33.800 ;
        RECT 115.800 33.100 116.200 33.200 ;
        RECT 116.700 33.100 117.000 34.900 ;
        RECT 118.200 34.800 119.400 34.900 ;
        RECT 117.400 34.100 117.800 34.600 ;
        RECT 118.200 34.100 118.600 34.200 ;
        RECT 117.400 33.800 118.600 34.100 ;
        RECT 119.800 33.100 120.200 39.900 ;
        RECT 122.700 36.200 123.100 39.900 ;
        RECT 123.400 36.800 123.800 37.200 ;
        RECT 123.500 36.200 123.800 36.800 ;
        RECT 122.700 35.900 123.200 36.200 ;
        RECT 123.500 35.900 124.200 36.200 ;
        RECT 124.600 35.900 125.000 39.900 ;
        RECT 125.400 36.200 125.800 39.900 ;
        RECT 127.000 36.200 127.400 39.900 ;
        RECT 127.800 37.900 128.200 39.900 ;
        RECT 127.900 37.800 128.200 37.900 ;
        RECT 129.400 37.900 129.800 39.900 ;
        RECT 131.800 37.900 132.200 39.900 ;
        RECT 129.400 37.800 129.700 37.900 ;
        RECT 127.900 37.500 129.700 37.800 ;
        RECT 131.900 37.800 132.200 37.900 ;
        RECT 133.400 37.900 133.800 39.900 ;
        RECT 133.400 37.800 133.700 37.900 ;
        RECT 131.900 37.500 133.700 37.800 ;
        RECT 127.900 36.200 128.200 37.500 ;
        RECT 128.600 37.100 129.000 37.200 ;
        RECT 132.600 37.100 133.000 37.200 ;
        RECT 128.600 36.800 133.000 37.100 ;
        RECT 128.600 36.400 129.000 36.800 ;
        RECT 132.600 36.400 133.000 36.800 ;
        RECT 133.400 36.200 133.700 37.500 ;
        RECT 125.400 35.900 127.400 36.200 ;
        RECT 122.200 34.400 122.600 35.200 ;
        RECT 122.900 34.200 123.200 35.900 ;
        RECT 123.800 35.800 124.200 35.900 ;
        RECT 124.700 35.200 125.000 35.900 ;
        RECT 127.800 35.800 128.200 36.200 ;
        RECT 126.600 35.200 127.000 35.400 ;
        RECT 124.600 34.900 125.800 35.200 ;
        RECT 126.600 35.100 127.400 35.200 ;
        RECT 127.900 35.100 128.200 35.800 ;
        RECT 130.200 35.400 130.600 36.200 ;
        RECT 131.000 35.400 131.400 36.200 ;
        RECT 133.400 35.800 133.800 36.200 ;
        RECT 134.200 35.900 134.600 39.900 ;
        RECT 135.000 36.200 135.400 39.900 ;
        RECT 136.600 36.200 137.000 39.900 ;
        RECT 137.400 37.900 137.800 39.900 ;
        RECT 137.500 37.800 137.800 37.900 ;
        RECT 139.000 37.900 139.400 39.900 ;
        RECT 139.000 37.800 139.300 37.900 ;
        RECT 137.500 37.500 139.300 37.800 ;
        RECT 137.500 36.200 137.800 37.500 ;
        RECT 138.200 36.400 138.600 37.200 ;
        RECT 140.600 36.200 141.000 39.900 ;
        RECT 142.200 36.200 142.600 39.900 ;
        RECT 135.000 35.900 137.000 36.200 ;
        RECT 133.400 35.200 133.700 35.800 ;
        RECT 134.300 35.200 134.600 35.900 ;
        RECT 137.400 35.800 137.800 36.200 ;
        RECT 139.000 36.100 139.400 36.200 ;
        RECT 139.800 36.100 140.200 36.200 ;
        RECT 139.000 35.800 140.200 36.100 ;
        RECT 140.600 35.900 142.600 36.200 ;
        RECT 143.000 35.900 143.400 39.900 ;
        RECT 144.600 37.900 145.000 39.900 ;
        RECT 144.700 37.800 145.000 37.900 ;
        RECT 146.200 37.900 146.600 39.900 ;
        RECT 146.200 37.800 146.500 37.900 ;
        RECT 144.700 37.500 146.500 37.800 ;
        RECT 145.400 36.400 145.800 37.200 ;
        RECT 146.200 36.200 146.500 37.500 ;
        RECT 147.400 36.800 147.800 37.200 ;
        RECT 147.400 36.200 147.700 36.800 ;
        RECT 148.100 36.200 148.500 39.900 ;
        RECT 136.200 35.200 136.600 35.400 ;
        RECT 126.600 34.900 128.200 35.100 ;
        RECT 124.600 34.800 125.000 34.900 ;
        RECT 120.600 33.400 121.000 34.200 ;
        RECT 121.400 34.100 121.800 34.200 ;
        RECT 122.900 34.100 124.200 34.200 ;
        RECT 124.600 34.100 125.000 34.200 ;
        RECT 121.400 33.800 122.200 34.100 ;
        RECT 122.900 33.800 125.000 34.100 ;
        RECT 121.800 33.600 122.200 33.800 ;
        RECT 121.500 33.100 123.300 33.300 ;
        RECT 123.800 33.100 124.100 33.800 ;
        RECT 112.600 33.000 114.600 33.100 ;
        RECT 112.600 31.100 113.000 33.000 ;
        RECT 114.200 31.100 114.600 33.000 ;
        RECT 115.000 32.800 116.200 33.100 ;
        RECT 115.000 31.100 115.400 32.800 ;
        RECT 115.900 32.400 116.300 32.800 ;
        RECT 116.600 31.100 117.000 33.100 ;
        RECT 119.300 32.800 120.200 33.100 ;
        RECT 121.400 33.000 123.400 33.100 ;
        RECT 119.300 32.200 119.700 32.800 ;
        RECT 119.000 31.800 119.700 32.200 ;
        RECT 119.300 31.100 119.700 31.800 ;
        RECT 121.400 31.100 121.800 33.000 ;
        RECT 123.000 31.100 123.400 33.000 ;
        RECT 123.800 31.100 124.200 33.100 ;
        RECT 124.600 32.800 125.000 33.200 ;
        RECT 125.500 33.100 125.800 34.900 ;
        RECT 127.000 34.800 128.200 34.900 ;
        RECT 128.600 34.800 129.800 35.200 ;
        RECT 131.800 34.800 132.600 35.200 ;
        RECT 133.400 34.800 133.800 35.200 ;
        RECT 134.200 34.900 135.400 35.200 ;
        RECT 136.200 34.900 137.000 35.200 ;
        RECT 134.200 34.800 134.600 34.900 ;
        RECT 126.200 33.800 126.600 34.600 ;
        RECT 127.900 34.200 128.200 34.800 ;
        RECT 133.400 34.200 133.700 34.800 ;
        RECT 127.900 34.100 128.700 34.200 ;
        RECT 132.900 34.100 133.700 34.200 ;
        RECT 127.900 33.900 128.800 34.100 ;
        RECT 124.700 32.400 125.100 32.800 ;
        RECT 125.400 31.100 125.800 33.100 ;
        RECT 128.400 31.100 128.800 33.900 ;
        RECT 132.800 33.900 133.700 34.100 ;
        RECT 134.200 34.100 134.600 34.200 ;
        RECT 135.100 34.100 135.400 34.900 ;
        RECT 136.600 34.800 137.000 34.900 ;
        RECT 132.800 33.100 133.200 33.900 ;
        RECT 134.200 33.800 135.400 34.100 ;
        RECT 135.800 33.800 136.200 34.600 ;
        RECT 137.500 34.200 137.800 35.800 ;
        RECT 139.800 35.400 140.200 35.800 ;
        RECT 141.000 35.200 141.400 35.400 ;
        RECT 143.000 35.200 143.300 35.900 ;
        RECT 143.800 35.400 144.200 36.200 ;
        RECT 146.200 35.800 146.600 36.200 ;
        RECT 147.000 35.900 147.700 36.200 ;
        RECT 148.000 35.900 148.500 36.200 ;
        RECT 147.000 35.800 147.400 35.900 ;
        RECT 138.600 34.800 139.400 35.200 ;
        RECT 140.600 34.900 141.400 35.200 ;
        RECT 142.200 34.900 143.400 35.200 ;
        RECT 140.600 34.800 141.000 34.900 ;
        RECT 137.500 34.100 138.300 34.200 ;
        RECT 137.500 33.900 139.300 34.100 ;
        RECT 138.000 33.800 139.300 33.900 ;
        RECT 141.400 33.800 141.800 34.600 ;
        RECT 134.200 33.100 134.600 33.200 ;
        RECT 135.100 33.100 135.400 33.800 ;
        RECT 132.800 32.800 134.600 33.100 ;
        RECT 132.800 31.100 133.200 32.800 ;
        RECT 134.300 32.400 134.700 32.800 ;
        RECT 135.000 31.100 135.400 33.100 ;
        RECT 138.000 31.100 138.400 33.800 ;
        RECT 139.000 33.200 139.300 33.800 ;
        RECT 139.000 32.800 139.400 33.200 ;
        RECT 142.200 33.100 142.500 34.900 ;
        RECT 143.000 34.800 143.400 34.900 ;
        RECT 144.600 34.800 145.400 35.200 ;
        RECT 143.000 34.200 143.300 34.800 ;
        RECT 146.200 34.200 146.500 35.800 ;
        RECT 148.000 34.200 148.300 35.900 ;
        RECT 148.600 34.400 149.000 35.200 ;
        RECT 143.000 33.800 143.400 34.200 ;
        RECT 145.700 34.100 146.500 34.200 ;
        RECT 145.600 33.900 146.500 34.100 ;
        RECT 142.200 31.100 142.600 33.100 ;
        RECT 143.000 32.800 143.400 33.200 ;
        RECT 142.900 32.400 143.300 32.800 ;
        RECT 145.600 32.200 146.000 33.900 ;
        RECT 147.000 33.800 148.300 34.200 ;
        RECT 149.400 34.100 149.800 34.200 ;
        RECT 150.200 34.100 150.600 34.200 ;
        RECT 149.000 33.800 150.600 34.100 ;
        RECT 147.100 33.100 147.400 33.800 ;
        RECT 149.000 33.600 149.400 33.800 ;
        RECT 147.900 33.100 149.700 33.300 ;
        RECT 145.400 31.800 146.000 32.200 ;
        RECT 145.600 31.100 146.000 31.800 ;
        RECT 147.000 31.100 147.400 33.100 ;
        RECT 147.800 33.000 149.800 33.100 ;
        RECT 147.800 31.100 148.200 33.000 ;
        RECT 149.400 31.100 149.800 33.000 ;
        RECT 1.400 27.600 1.800 29.900 ;
        RECT 3.000 27.600 3.400 29.900 ;
        RECT 4.600 27.600 5.000 29.900 ;
        RECT 6.200 27.600 6.600 29.900 ;
        RECT 7.800 27.900 8.200 29.900 ;
        RECT 10.000 28.100 10.800 29.900 ;
        RECT 7.800 27.600 9.000 27.900 ;
        RECT 1.400 27.200 2.300 27.600 ;
        RECT 3.000 27.200 4.100 27.600 ;
        RECT 4.600 27.200 5.700 27.600 ;
        RECT 6.200 27.200 7.400 27.600 ;
        RECT 8.600 27.500 9.000 27.600 ;
        RECT 9.300 27.400 9.700 27.800 ;
        RECT 9.300 27.200 9.600 27.400 ;
        RECT 1.900 26.900 2.300 27.200 ;
        RECT 3.700 26.900 4.100 27.200 ;
        RECT 5.300 26.900 5.700 27.200 ;
        RECT 1.900 26.500 3.200 26.900 ;
        RECT 3.700 26.500 4.900 26.900 ;
        RECT 5.300 26.500 6.600 26.900 ;
        RECT 1.900 25.800 2.300 26.500 ;
        RECT 3.700 25.800 4.100 26.500 ;
        RECT 5.300 25.800 5.700 26.500 ;
        RECT 7.000 25.800 7.400 27.200 ;
        RECT 7.800 26.800 8.600 27.200 ;
        RECT 9.200 26.800 9.600 27.200 ;
        RECT 10.000 26.400 10.300 28.100 ;
        RECT 12.600 27.900 13.000 29.900 ;
        RECT 10.600 27.700 11.400 27.800 ;
        RECT 10.600 27.400 11.600 27.700 ;
        RECT 11.900 27.600 13.000 27.900 ;
        RECT 11.900 27.500 12.300 27.600 ;
        RECT 13.400 27.500 13.800 29.900 ;
        RECT 15.600 29.200 16.000 29.900 ;
        RECT 15.000 28.900 16.000 29.200 ;
        RECT 17.800 28.900 18.200 29.900 ;
        RECT 19.900 29.200 20.500 29.900 ;
        RECT 19.800 28.900 20.500 29.200 ;
        RECT 15.000 28.500 15.400 28.900 ;
        RECT 17.800 28.600 18.100 28.900 ;
        RECT 15.800 28.200 16.200 28.600 ;
        RECT 16.700 28.300 18.100 28.600 ;
        RECT 19.800 28.500 20.200 28.900 ;
        RECT 16.700 28.200 17.100 28.300 ;
        RECT 11.300 27.200 11.600 27.400 ;
        RECT 10.600 26.700 11.000 27.100 ;
        RECT 11.300 26.900 13.000 27.200 ;
        RECT 12.200 26.800 13.000 26.900 ;
        RECT 13.800 27.100 14.600 27.200 ;
        RECT 15.900 27.100 16.200 28.200 ;
        RECT 20.700 27.700 21.100 27.800 ;
        RECT 22.200 27.700 22.600 29.900 ;
        RECT 20.700 27.400 22.600 27.700 ;
        RECT 23.000 27.500 23.400 29.900 ;
        RECT 25.200 29.200 25.600 29.900 ;
        RECT 24.600 28.900 25.600 29.200 ;
        RECT 27.400 28.900 27.800 29.900 ;
        RECT 29.500 29.200 30.100 29.900 ;
        RECT 29.400 28.900 30.100 29.200 ;
        RECT 24.600 28.500 25.000 28.900 ;
        RECT 27.400 28.600 27.700 28.900 ;
        RECT 25.400 28.200 25.800 28.600 ;
        RECT 26.300 28.300 27.700 28.600 ;
        RECT 29.400 28.500 29.800 28.900 ;
        RECT 26.300 28.200 26.700 28.300 ;
        RECT 18.700 27.100 19.100 27.200 ;
        RECT 13.800 26.800 19.300 27.100 ;
        RECT 15.300 26.700 15.700 26.800 ;
        RECT 9.800 26.200 10.300 26.400 ;
        RECT 9.400 26.100 10.300 26.200 ;
        RECT 10.700 26.400 11.000 26.700 ;
        RECT 10.700 26.100 12.000 26.400 ;
        RECT 9.400 25.800 10.100 26.100 ;
        RECT 11.600 26.000 12.000 26.100 ;
        RECT 14.500 26.200 14.900 26.300 ;
        RECT 15.800 26.200 16.200 26.300 ;
        RECT 14.500 25.900 17.000 26.200 ;
        RECT 16.600 25.800 17.000 25.900 ;
        RECT 1.400 25.400 2.300 25.800 ;
        RECT 3.000 25.400 4.100 25.800 ;
        RECT 4.600 25.400 5.700 25.800 ;
        RECT 6.200 25.400 7.400 25.800 ;
        RECT 1.400 21.100 1.800 25.400 ;
        RECT 3.000 21.100 3.400 25.400 ;
        RECT 4.600 21.100 5.000 25.400 ;
        RECT 6.200 21.100 6.600 25.400 ;
        RECT 9.800 25.100 10.100 25.800 ;
        RECT 10.500 25.700 10.900 25.800 ;
        RECT 10.500 25.400 12.200 25.700 ;
        RECT 11.900 25.100 12.200 25.400 ;
        RECT 13.400 25.500 16.200 25.600 ;
        RECT 13.400 25.400 16.300 25.500 ;
        RECT 13.400 25.300 18.300 25.400 ;
        RECT 7.800 24.800 9.000 25.100 ;
        RECT 9.800 24.800 10.800 25.100 ;
        RECT 7.800 21.100 8.200 24.800 ;
        RECT 8.600 24.700 9.000 24.800 ;
        RECT 10.000 21.100 10.800 24.800 ;
        RECT 11.900 24.800 13.000 25.100 ;
        RECT 11.900 24.700 12.300 24.800 ;
        RECT 12.600 21.100 13.000 24.800 ;
        RECT 13.400 21.100 13.800 25.300 ;
        RECT 15.900 25.100 18.300 25.300 ;
        RECT 15.000 24.500 17.700 24.800 ;
        RECT 15.000 24.400 15.400 24.500 ;
        RECT 17.300 24.400 17.700 24.500 ;
        RECT 18.000 24.500 18.300 25.100 ;
        RECT 19.000 25.200 19.300 26.800 ;
        RECT 19.800 26.400 20.200 26.500 ;
        RECT 19.800 26.100 21.700 26.400 ;
        RECT 21.300 26.000 21.700 26.100 ;
        RECT 20.500 25.700 20.900 25.800 ;
        RECT 22.200 25.700 22.600 27.400 ;
        RECT 23.400 27.100 24.200 27.200 ;
        RECT 25.500 27.100 25.800 28.200 ;
        RECT 30.300 27.700 30.700 27.800 ;
        RECT 31.800 27.700 32.200 29.900 ;
        RECT 30.300 27.400 32.200 27.700 ;
        RECT 32.600 27.500 33.000 29.900 ;
        RECT 34.800 29.200 35.200 29.900 ;
        RECT 34.200 28.900 35.200 29.200 ;
        RECT 37.000 28.900 37.400 29.900 ;
        RECT 39.100 29.200 39.700 29.900 ;
        RECT 39.000 28.900 39.700 29.200 ;
        RECT 34.200 28.500 34.600 28.900 ;
        RECT 37.000 28.600 37.300 28.900 ;
        RECT 35.000 28.200 35.400 28.600 ;
        RECT 35.900 28.300 37.300 28.600 ;
        RECT 39.000 28.500 39.400 28.900 ;
        RECT 35.900 28.200 36.300 28.300 ;
        RECT 28.300 27.100 28.700 27.200 ;
        RECT 23.400 26.800 28.900 27.100 ;
        RECT 24.900 26.700 25.300 26.800 ;
        RECT 24.100 26.200 24.500 26.300 ;
        RECT 25.400 26.200 25.800 26.300 ;
        RECT 24.100 25.900 26.600 26.200 ;
        RECT 26.200 25.800 26.600 25.900 ;
        RECT 20.500 25.400 22.600 25.700 ;
        RECT 19.000 24.900 20.200 25.200 ;
        RECT 18.700 24.500 19.100 24.600 ;
        RECT 18.000 24.200 19.100 24.500 ;
        RECT 19.900 24.400 20.200 24.900 ;
        RECT 19.900 24.200 20.600 24.400 ;
        RECT 19.900 24.000 21.000 24.200 ;
        RECT 20.300 23.800 21.000 24.000 ;
        RECT 16.700 23.700 17.100 23.800 ;
        RECT 18.100 23.700 18.500 23.800 ;
        RECT 15.000 23.100 15.400 23.500 ;
        RECT 16.700 23.400 18.500 23.700 ;
        RECT 17.800 23.100 18.100 23.400 ;
        RECT 19.800 23.100 20.200 23.500 ;
        RECT 15.000 22.800 16.000 23.100 ;
        RECT 15.600 21.100 16.000 22.800 ;
        RECT 17.800 21.100 18.200 23.100 ;
        RECT 19.900 21.100 20.500 23.100 ;
        RECT 22.200 21.100 22.600 25.400 ;
        RECT 23.000 25.500 25.800 25.600 ;
        RECT 23.000 25.400 25.900 25.500 ;
        RECT 23.000 25.300 27.900 25.400 ;
        RECT 23.000 21.100 23.400 25.300 ;
        RECT 25.500 25.100 27.900 25.300 ;
        RECT 24.600 24.500 27.300 24.800 ;
        RECT 24.600 24.400 25.000 24.500 ;
        RECT 26.900 24.400 27.300 24.500 ;
        RECT 27.600 24.500 27.900 25.100 ;
        RECT 28.600 25.200 28.900 26.800 ;
        RECT 29.400 26.400 29.800 26.500 ;
        RECT 29.400 26.100 31.300 26.400 ;
        RECT 30.900 26.000 31.300 26.100 ;
        RECT 30.100 25.700 30.500 25.800 ;
        RECT 31.800 25.700 32.200 27.400 ;
        RECT 33.000 27.100 33.800 27.200 ;
        RECT 35.100 27.100 35.400 28.200 ;
        RECT 39.900 27.700 40.300 27.800 ;
        RECT 41.400 27.700 41.800 29.900 ;
        RECT 39.900 27.400 41.800 27.700 ;
        RECT 42.200 27.500 42.600 29.900 ;
        RECT 44.400 29.200 44.800 29.900 ;
        RECT 43.800 28.900 44.800 29.200 ;
        RECT 46.600 28.900 47.000 29.900 ;
        RECT 48.700 29.200 49.300 29.900 ;
        RECT 48.600 28.900 49.300 29.200 ;
        RECT 43.800 28.500 44.200 28.900 ;
        RECT 46.600 28.600 46.900 28.900 ;
        RECT 44.600 28.200 45.000 28.600 ;
        RECT 45.500 28.300 46.900 28.600 ;
        RECT 48.600 28.500 49.000 28.900 ;
        RECT 45.500 28.200 45.900 28.300 ;
        RECT 37.900 27.100 38.300 27.200 ;
        RECT 33.000 26.800 38.500 27.100 ;
        RECT 34.500 26.700 34.900 26.800 ;
        RECT 33.700 26.200 34.100 26.300 ;
        RECT 35.000 26.200 35.400 26.300 ;
        RECT 33.700 25.900 36.200 26.200 ;
        RECT 35.800 25.800 36.200 25.900 ;
        RECT 30.100 25.400 32.200 25.700 ;
        RECT 28.600 24.900 29.800 25.200 ;
        RECT 28.300 24.500 28.700 24.600 ;
        RECT 27.600 24.200 28.700 24.500 ;
        RECT 29.500 24.400 29.800 24.900 ;
        RECT 29.500 24.000 30.200 24.400 ;
        RECT 26.300 23.700 26.700 23.800 ;
        RECT 27.700 23.700 28.100 23.800 ;
        RECT 24.600 23.100 25.000 23.500 ;
        RECT 26.300 23.400 28.100 23.700 ;
        RECT 27.400 23.100 27.700 23.400 ;
        RECT 29.400 23.100 29.800 23.500 ;
        RECT 24.600 22.800 25.600 23.100 ;
        RECT 25.200 21.100 25.600 22.800 ;
        RECT 27.400 21.100 27.800 23.100 ;
        RECT 29.500 21.100 30.100 23.100 ;
        RECT 31.800 21.100 32.200 25.400 ;
        RECT 32.600 25.500 35.400 25.600 ;
        RECT 32.600 25.400 35.500 25.500 ;
        RECT 32.600 25.300 37.500 25.400 ;
        RECT 32.600 21.100 33.000 25.300 ;
        RECT 35.100 25.100 37.500 25.300 ;
        RECT 34.200 24.500 36.900 24.800 ;
        RECT 34.200 24.400 34.600 24.500 ;
        RECT 36.500 24.400 36.900 24.500 ;
        RECT 37.200 24.500 37.500 25.100 ;
        RECT 38.200 25.200 38.500 26.800 ;
        RECT 39.000 26.400 39.400 26.500 ;
        RECT 39.000 26.100 40.900 26.400 ;
        RECT 40.500 26.000 40.900 26.100 ;
        RECT 39.700 25.700 40.100 25.800 ;
        RECT 41.400 25.700 41.800 27.400 ;
        RECT 42.600 27.100 43.400 27.200 ;
        RECT 44.700 27.100 45.000 28.200 ;
        RECT 49.500 27.700 49.900 27.800 ;
        RECT 51.000 27.700 51.400 29.900 ;
        RECT 49.500 27.400 51.400 27.700 ;
        RECT 53.400 27.500 53.800 29.900 ;
        RECT 55.600 29.200 56.000 29.900 ;
        RECT 55.000 28.900 56.000 29.200 ;
        RECT 57.800 28.900 58.200 29.900 ;
        RECT 59.900 29.200 60.500 29.900 ;
        RECT 59.800 28.900 60.500 29.200 ;
        RECT 55.000 28.500 55.400 28.900 ;
        RECT 57.800 28.600 58.100 28.900 ;
        RECT 55.800 28.200 56.200 28.600 ;
        RECT 56.700 28.300 58.100 28.600 ;
        RECT 59.800 28.500 60.200 28.900 ;
        RECT 56.700 28.200 57.100 28.300 ;
        RECT 47.500 27.100 47.900 27.200 ;
        RECT 42.600 26.800 48.100 27.100 ;
        RECT 44.100 26.700 44.500 26.800 ;
        RECT 43.300 26.200 43.700 26.300 ;
        RECT 44.600 26.200 45.000 26.300 ;
        RECT 47.800 26.200 48.100 26.800 ;
        RECT 48.600 26.400 49.000 26.500 ;
        RECT 43.300 25.900 45.800 26.200 ;
        RECT 45.400 25.800 45.800 25.900 ;
        RECT 47.800 25.800 48.200 26.200 ;
        RECT 48.600 26.100 50.500 26.400 ;
        RECT 50.100 26.000 50.500 26.100 ;
        RECT 39.700 25.400 41.800 25.700 ;
        RECT 38.200 24.900 39.400 25.200 ;
        RECT 37.900 24.500 38.300 24.600 ;
        RECT 37.200 24.200 38.300 24.500 ;
        RECT 39.100 24.400 39.400 24.900 ;
        RECT 39.100 24.000 39.800 24.400 ;
        RECT 35.900 23.700 36.300 23.800 ;
        RECT 37.300 23.700 37.700 23.800 ;
        RECT 34.200 23.100 34.600 23.500 ;
        RECT 35.900 23.400 37.700 23.700 ;
        RECT 37.000 23.100 37.300 23.400 ;
        RECT 39.000 23.100 39.400 23.500 ;
        RECT 34.200 22.800 35.200 23.100 ;
        RECT 34.800 21.100 35.200 22.800 ;
        RECT 37.000 21.100 37.400 23.100 ;
        RECT 39.100 21.100 39.700 23.100 ;
        RECT 41.400 21.100 41.800 25.400 ;
        RECT 42.200 25.500 45.000 25.600 ;
        RECT 42.200 25.400 45.100 25.500 ;
        RECT 42.200 25.300 47.100 25.400 ;
        RECT 42.200 21.100 42.600 25.300 ;
        RECT 44.700 25.100 47.100 25.300 ;
        RECT 43.800 24.500 46.500 24.800 ;
        RECT 43.800 24.400 44.200 24.500 ;
        RECT 46.100 24.400 46.500 24.500 ;
        RECT 46.800 24.500 47.100 25.100 ;
        RECT 47.800 25.200 48.100 25.800 ;
        RECT 49.300 25.700 49.700 25.800 ;
        RECT 51.000 25.700 51.400 27.400 ;
        RECT 53.800 27.100 54.600 27.200 ;
        RECT 55.900 27.100 56.200 28.200 ;
        RECT 60.700 27.700 61.100 27.800 ;
        RECT 62.200 27.700 62.600 29.900 ;
        RECT 60.700 27.400 62.600 27.700 ;
        RECT 63.800 27.600 64.200 29.900 ;
        RECT 65.400 27.600 65.800 29.900 ;
        RECT 67.000 27.600 67.400 29.900 ;
        RECT 68.600 27.600 69.000 29.900 ;
        RECT 57.400 27.100 57.800 27.200 ;
        RECT 58.700 27.100 59.100 27.200 ;
        RECT 53.800 26.800 59.300 27.100 ;
        RECT 55.300 26.700 55.700 26.800 ;
        RECT 54.500 26.200 54.900 26.300 ;
        RECT 55.800 26.200 56.200 26.300 ;
        RECT 54.500 25.900 57.000 26.200 ;
        RECT 56.600 25.800 57.000 25.900 ;
        RECT 49.300 25.400 51.400 25.700 ;
        RECT 47.800 24.900 49.000 25.200 ;
        RECT 47.500 24.500 47.900 24.600 ;
        RECT 46.800 24.200 47.900 24.500 ;
        RECT 48.700 24.400 49.000 24.900 ;
        RECT 48.700 24.000 49.400 24.400 ;
        RECT 45.500 23.700 45.900 23.800 ;
        RECT 46.900 23.700 47.300 23.800 ;
        RECT 43.800 23.100 44.200 23.500 ;
        RECT 45.500 23.400 47.300 23.700 ;
        RECT 46.600 23.100 46.900 23.400 ;
        RECT 48.600 23.100 49.000 23.500 ;
        RECT 43.800 22.800 44.800 23.100 ;
        RECT 44.400 21.100 44.800 22.800 ;
        RECT 46.600 21.100 47.000 23.100 ;
        RECT 48.700 21.100 49.300 23.100 ;
        RECT 51.000 21.100 51.400 25.400 ;
        RECT 53.400 25.500 56.200 25.600 ;
        RECT 53.400 25.400 56.300 25.500 ;
        RECT 53.400 25.300 58.300 25.400 ;
        RECT 53.400 21.100 53.800 25.300 ;
        RECT 55.900 25.100 58.300 25.300 ;
        RECT 55.000 24.500 57.700 24.800 ;
        RECT 55.000 24.400 55.400 24.500 ;
        RECT 57.300 24.400 57.700 24.500 ;
        RECT 58.000 24.500 58.300 25.100 ;
        RECT 59.000 25.200 59.300 26.800 ;
        RECT 59.800 26.400 60.200 26.500 ;
        RECT 59.800 26.100 61.700 26.400 ;
        RECT 61.300 26.000 61.700 26.100 ;
        RECT 60.500 25.700 60.900 25.800 ;
        RECT 62.200 25.700 62.600 27.400 ;
        RECT 60.500 25.400 62.600 25.700 ;
        RECT 63.000 27.200 64.200 27.600 ;
        RECT 64.700 27.200 65.800 27.600 ;
        RECT 66.300 27.200 67.400 27.600 ;
        RECT 68.100 27.200 69.000 27.600 ;
        RECT 71.000 27.600 71.400 29.900 ;
        RECT 72.600 27.600 73.000 29.900 ;
        RECT 74.200 27.600 74.600 29.900 ;
        RECT 75.800 27.600 76.200 29.900 ;
        RECT 77.400 27.900 77.800 29.900 ;
        RECT 79.600 28.100 80.400 29.900 ;
        RECT 77.400 27.600 78.500 27.900 ;
        RECT 79.000 27.700 79.800 27.800 ;
        RECT 71.000 27.200 71.900 27.600 ;
        RECT 72.600 27.200 73.700 27.600 ;
        RECT 74.200 27.200 75.300 27.600 ;
        RECT 75.800 27.200 77.000 27.600 ;
        RECT 78.100 27.500 78.500 27.600 ;
        RECT 78.800 27.400 79.800 27.700 ;
        RECT 78.800 27.200 79.100 27.400 ;
        RECT 63.000 25.800 63.400 27.200 ;
        RECT 64.700 26.900 65.100 27.200 ;
        RECT 66.300 26.900 66.700 27.200 ;
        RECT 68.100 26.900 68.500 27.200 ;
        RECT 63.800 26.500 65.100 26.900 ;
        RECT 65.500 26.500 66.700 26.900 ;
        RECT 67.200 26.500 68.500 26.900 ;
        RECT 64.700 25.800 65.100 26.500 ;
        RECT 66.300 25.800 66.700 26.500 ;
        RECT 68.100 25.800 68.500 26.500 ;
        RECT 71.500 26.900 71.900 27.200 ;
        RECT 73.300 26.900 73.700 27.200 ;
        RECT 74.900 26.900 75.300 27.200 ;
        RECT 71.500 26.500 72.800 26.900 ;
        RECT 73.300 26.500 74.500 26.900 ;
        RECT 74.900 26.500 76.200 26.900 ;
        RECT 71.500 25.800 71.900 26.500 ;
        RECT 73.300 25.800 73.700 26.500 ;
        RECT 74.900 25.800 75.300 26.500 ;
        RECT 76.600 25.800 77.000 27.200 ;
        RECT 77.400 26.900 79.100 27.200 ;
        RECT 77.400 26.800 78.200 26.900 ;
        RECT 79.400 26.700 79.800 27.100 ;
        RECT 79.400 26.400 79.700 26.700 ;
        RECT 78.400 26.100 79.700 26.400 ;
        RECT 80.100 26.400 80.400 28.100 ;
        RECT 82.200 27.900 82.600 29.900 ;
        RECT 80.700 27.400 81.100 27.800 ;
        RECT 81.400 27.600 82.600 27.900 ;
        RECT 81.400 27.500 81.800 27.600 ;
        RECT 80.800 27.200 81.100 27.400 ;
        RECT 80.800 26.800 81.200 27.200 ;
        RECT 81.800 27.100 82.600 27.200 ;
        RECT 83.000 27.100 83.400 29.900 ;
        RECT 83.800 27.800 84.200 28.600 ;
        RECT 84.700 28.200 85.100 28.600 ;
        RECT 84.600 27.800 85.000 28.200 ;
        RECT 85.400 27.800 85.800 29.900 ;
        RECT 81.800 26.800 83.400 27.100 ;
        RECT 80.100 26.200 80.600 26.400 ;
        RECT 80.100 26.100 81.000 26.200 ;
        RECT 78.400 26.000 78.800 26.100 ;
        RECT 80.300 25.800 81.000 26.100 ;
        RECT 63.000 25.400 64.200 25.800 ;
        RECT 64.700 25.400 65.800 25.800 ;
        RECT 66.300 25.400 67.400 25.800 ;
        RECT 68.100 25.400 69.000 25.800 ;
        RECT 59.000 24.900 60.200 25.200 ;
        RECT 58.700 24.500 59.100 24.600 ;
        RECT 58.000 24.200 59.100 24.500 ;
        RECT 59.900 24.400 60.200 24.900 ;
        RECT 59.900 24.000 60.600 24.400 ;
        RECT 56.700 23.700 57.100 23.800 ;
        RECT 58.100 23.700 58.500 23.800 ;
        RECT 55.000 23.100 55.400 23.500 ;
        RECT 56.700 23.400 58.500 23.700 ;
        RECT 57.800 23.100 58.100 23.400 ;
        RECT 59.800 23.100 60.200 23.500 ;
        RECT 55.000 22.800 56.000 23.100 ;
        RECT 55.600 21.100 56.000 22.800 ;
        RECT 57.800 21.100 58.200 23.100 ;
        RECT 59.900 21.100 60.500 23.100 ;
        RECT 62.200 21.100 62.600 25.400 ;
        RECT 63.800 21.100 64.200 25.400 ;
        RECT 65.400 21.100 65.800 25.400 ;
        RECT 67.000 21.100 67.400 25.400 ;
        RECT 68.600 21.100 69.000 25.400 ;
        RECT 71.000 25.400 71.900 25.800 ;
        RECT 72.600 25.400 73.700 25.800 ;
        RECT 74.200 25.400 75.300 25.800 ;
        RECT 75.800 25.400 77.000 25.800 ;
        RECT 79.500 25.700 79.900 25.800 ;
        RECT 78.200 25.400 79.900 25.700 ;
        RECT 71.000 21.100 71.400 25.400 ;
        RECT 72.600 21.100 73.000 25.400 ;
        RECT 74.200 21.100 74.600 25.400 ;
        RECT 75.800 21.100 76.200 25.400 ;
        RECT 78.200 25.100 78.500 25.400 ;
        RECT 80.300 25.100 80.600 25.800 ;
        RECT 77.400 24.800 78.500 25.100 ;
        RECT 77.400 21.100 77.800 24.800 ;
        RECT 78.100 24.700 78.500 24.800 ;
        RECT 79.600 24.800 80.600 25.100 ;
        RECT 81.400 24.800 82.600 25.100 ;
        RECT 79.600 21.100 80.400 24.800 ;
        RECT 81.400 24.700 81.800 24.800 ;
        RECT 82.200 21.100 82.600 24.800 ;
        RECT 83.000 21.100 83.400 26.800 ;
        RECT 84.600 26.100 85.000 26.200 ;
        RECT 85.500 26.100 85.800 27.800 ;
        RECT 88.600 28.900 89.000 29.900 ;
        RECT 88.600 27.200 88.900 28.900 ;
        RECT 89.400 27.800 89.800 28.600 ;
        RECT 90.200 27.800 90.600 28.600 ;
        RECT 86.200 26.400 86.600 27.200 ;
        RECT 88.600 27.100 89.000 27.200 ;
        RECT 87.000 26.800 89.000 27.100 ;
        RECT 89.400 27.100 89.700 27.800 ;
        RECT 91.000 27.100 91.400 29.900 ;
        RECT 91.800 27.900 92.200 29.900 ;
        RECT 92.600 28.000 93.000 29.900 ;
        RECT 94.200 28.000 94.600 29.900 ;
        RECT 95.100 28.200 95.500 28.600 ;
        RECT 92.600 27.900 94.600 28.000 ;
        RECT 91.900 27.200 92.200 27.900 ;
        RECT 92.700 27.700 94.500 27.900 ;
        RECT 95.000 27.800 95.400 28.200 ;
        RECT 95.800 27.900 96.200 29.900 ;
        RECT 93.800 27.200 94.200 27.400 ;
        RECT 95.900 27.200 96.200 27.900 ;
        RECT 89.400 26.800 91.400 27.100 ;
        RECT 91.800 26.800 93.100 27.200 ;
        RECT 93.800 27.100 94.600 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 93.800 26.900 96.200 27.100 ;
        RECT 94.200 26.800 96.200 26.900 ;
        RECT 87.000 26.200 87.300 26.800 ;
        RECT 87.000 26.100 87.400 26.200 ;
        RECT 84.600 25.800 85.800 26.100 ;
        RECT 86.600 25.800 87.400 26.100 ;
        RECT 84.700 25.100 85.000 25.800 ;
        RECT 86.600 25.600 87.000 25.800 ;
        RECT 87.800 25.400 88.200 26.200 ;
        RECT 88.600 25.100 88.900 26.800 ;
        RECT 84.600 21.100 85.000 25.100 ;
        RECT 85.400 24.800 87.400 25.100 ;
        RECT 85.400 21.100 85.800 24.800 ;
        RECT 87.000 21.100 87.400 24.800 ;
        RECT 88.100 24.700 89.000 25.100 ;
        RECT 88.100 21.100 88.500 24.700 ;
        RECT 91.000 21.100 91.400 26.800 ;
        RECT 92.800 26.200 93.100 26.800 ;
        RECT 92.600 25.800 93.100 26.200 ;
        RECT 93.400 25.800 93.800 26.600 ;
        RECT 95.000 26.100 95.400 26.200 ;
        RECT 95.900 26.100 96.200 26.800 ;
        RECT 96.600 27.100 97.000 27.200 ;
        RECT 97.400 27.100 97.800 27.200 ;
        RECT 98.800 27.100 99.200 29.900 ;
        RECT 103.100 28.200 103.500 28.600 ;
        RECT 103.000 27.800 103.400 28.200 ;
        RECT 103.800 27.900 104.200 29.900 ;
        RECT 96.600 26.800 97.800 27.100 ;
        RECT 98.300 26.900 99.200 27.100 ;
        RECT 98.300 26.800 99.100 26.900 ;
        RECT 96.600 26.400 97.000 26.800 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 95.000 25.800 96.200 26.100 ;
        RECT 97.000 25.800 97.800 26.100 ;
        RECT 91.800 25.100 92.200 25.200 ;
        RECT 92.800 25.100 93.100 25.800 ;
        RECT 95.100 25.100 95.400 25.800 ;
        RECT 97.000 25.600 97.400 25.800 ;
        RECT 98.300 25.200 98.600 26.800 ;
        RECT 99.400 25.800 100.200 26.200 ;
        RECT 103.000 26.100 103.400 26.200 ;
        RECT 103.900 26.100 104.200 27.900 ;
        RECT 104.600 26.400 105.000 27.200 ;
        RECT 106.800 27.100 107.200 29.900 ;
        RECT 106.300 26.900 107.200 27.100 ;
        RECT 106.300 26.800 107.100 26.900 ;
        RECT 105.400 26.100 105.800 26.200 ;
        RECT 103.000 25.800 104.200 26.100 ;
        RECT 105.000 25.800 105.800 26.100 ;
        RECT 91.800 24.800 92.500 25.100 ;
        RECT 92.800 24.800 93.300 25.100 ;
        RECT 92.200 24.200 92.500 24.800 ;
        RECT 92.200 23.800 92.600 24.200 ;
        RECT 92.900 21.100 93.300 24.800 ;
        RECT 95.000 21.100 95.400 25.100 ;
        RECT 95.800 24.800 97.800 25.100 ;
        RECT 98.200 24.800 98.600 25.200 ;
        RECT 100.600 24.800 101.000 25.600 ;
        RECT 103.100 25.100 103.400 25.800 ;
        RECT 105.000 25.600 105.400 25.800 ;
        RECT 106.300 25.200 106.600 26.800 ;
        RECT 107.400 25.800 108.200 26.200 ;
        RECT 95.800 21.100 96.200 24.800 ;
        RECT 97.400 21.100 97.800 24.800 ;
        RECT 98.300 23.500 98.600 24.800 ;
        RECT 99.000 23.800 99.400 24.600 ;
        RECT 98.300 23.200 100.100 23.500 ;
        RECT 98.300 23.100 98.600 23.200 ;
        RECT 98.200 21.100 98.600 23.100 ;
        RECT 99.800 21.100 100.200 23.200 ;
        RECT 103.000 21.100 103.400 25.100 ;
        RECT 103.800 24.800 105.800 25.100 ;
        RECT 106.200 24.800 106.600 25.200 ;
        RECT 108.600 25.100 109.000 26.200 ;
        RECT 109.400 25.100 109.800 29.900 ;
        RECT 111.800 28.900 112.200 29.900 ;
        RECT 114.200 28.900 114.600 29.900 ;
        RECT 110.200 27.800 110.600 28.600 ;
        RECT 111.000 27.800 111.400 28.600 ;
        RECT 111.900 27.200 112.200 28.900 ;
        RECT 113.400 27.800 113.800 28.600 ;
        RECT 114.300 27.800 114.600 28.900 ;
        RECT 115.800 27.900 116.200 29.900 ;
        RECT 119.000 28.900 119.400 29.900 ;
        RECT 120.600 29.200 121.000 29.900 ;
        RECT 114.300 27.500 115.500 27.800 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 114.200 26.800 114.700 27.200 ;
        RECT 110.200 26.100 110.600 26.200 ;
        RECT 111.900 26.100 112.200 26.800 ;
        RECT 114.400 26.400 114.800 26.800 ;
        RECT 110.200 25.800 112.200 26.100 ;
        RECT 111.900 25.100 112.200 25.800 ;
        RECT 112.600 25.400 113.000 26.200 ;
        RECT 115.200 26.000 115.500 27.500 ;
        RECT 115.900 27.100 116.200 27.900 ;
        RECT 118.800 28.800 119.400 28.900 ;
        RECT 120.500 28.900 121.000 29.200 ;
        RECT 120.500 28.800 120.800 28.900 ;
        RECT 118.800 28.500 120.800 28.800 ;
        RECT 118.800 27.200 119.100 28.500 ;
        RECT 120.900 27.800 121.800 28.200 ;
        RECT 123.000 28.000 123.400 29.900 ;
        RECT 124.600 28.000 125.000 29.900 ;
        RECT 123.000 27.900 125.000 28.000 ;
        RECT 125.400 27.900 125.800 29.900 ;
        RECT 127.000 28.900 127.400 29.900 ;
        RECT 116.600 27.100 117.000 27.200 ;
        RECT 115.800 26.800 117.000 27.100 ;
        RECT 118.800 26.800 119.400 27.200 ;
        RECT 120.200 26.800 121.000 27.200 ;
        RECT 121.400 27.100 121.700 27.800 ;
        RECT 123.100 27.700 124.900 27.900 ;
        RECT 123.400 27.200 123.800 27.400 ;
        RECT 125.400 27.200 125.700 27.900 ;
        RECT 126.200 27.800 126.600 28.600 ;
        RECT 127.100 27.200 127.400 28.900 ;
        RECT 130.100 27.900 130.900 29.900 ;
        RECT 133.400 28.900 133.800 29.900 ;
        RECT 123.000 27.100 123.800 27.200 ;
        RECT 121.400 26.900 123.800 27.100 ;
        RECT 121.400 26.800 123.400 26.900 ;
        RECT 124.500 26.800 125.800 27.200 ;
        RECT 127.000 27.100 127.400 27.200 ;
        RECT 127.000 26.800 128.900 27.100 ;
        RECT 115.900 26.200 116.200 26.800 ;
        RECT 115.100 25.700 115.500 26.000 ;
        RECT 115.800 25.800 116.200 26.200 ;
        RECT 113.400 25.600 115.500 25.700 ;
        RECT 113.400 25.400 115.400 25.600 ;
        RECT 108.600 24.800 109.800 25.100 ;
        RECT 103.800 21.100 104.200 24.800 ;
        RECT 105.400 21.100 105.800 24.800 ;
        RECT 106.300 23.500 106.600 24.800 ;
        RECT 107.000 23.800 107.400 24.600 ;
        RECT 106.300 23.200 108.100 23.500 ;
        RECT 106.300 23.100 106.600 23.200 ;
        RECT 106.200 21.100 106.600 23.100 ;
        RECT 107.800 23.100 108.100 23.200 ;
        RECT 107.800 21.100 108.200 23.100 ;
        RECT 109.400 21.100 109.800 24.800 ;
        RECT 111.800 24.700 112.700 25.100 ;
        RECT 112.300 21.100 112.700 24.700 ;
        RECT 113.400 21.100 113.800 25.400 ;
        RECT 115.900 25.100 116.200 25.800 ;
        RECT 118.800 25.200 119.100 26.800 ;
        RECT 119.400 26.100 120.200 26.200 ;
        RECT 123.000 26.100 123.400 26.200 ;
        RECT 123.800 26.100 124.200 26.600 ;
        RECT 119.400 25.800 124.200 26.100 ;
        RECT 124.500 26.100 124.800 26.800 ;
        RECT 126.200 26.100 126.600 26.200 ;
        RECT 124.500 25.800 126.600 26.100 ;
        RECT 115.500 24.800 116.200 25.100 ;
        RECT 117.400 24.900 119.100 25.200 ;
        RECT 124.500 25.100 124.800 25.800 ;
        RECT 125.400 25.100 125.800 25.200 ;
        RECT 127.100 25.100 127.400 26.800 ;
        RECT 128.600 26.200 128.900 26.800 ;
        RECT 129.400 26.400 129.800 27.200 ;
        RECT 130.300 26.200 130.600 27.900 ;
        RECT 133.400 27.200 133.700 28.900 ;
        RECT 134.200 27.800 134.600 28.600 ;
        RECT 131.000 26.800 131.400 27.200 ;
        RECT 133.400 26.800 133.800 27.200 ;
        RECT 135.600 27.100 136.000 29.900 ;
        RECT 138.200 28.000 138.600 29.900 ;
        RECT 139.800 28.000 140.200 29.900 ;
        RECT 138.200 27.900 140.200 28.000 ;
        RECT 140.600 27.900 141.000 29.900 ;
        RECT 141.700 28.200 142.100 29.900 ;
        RECT 141.700 27.900 142.600 28.200 ;
        RECT 138.300 27.700 140.100 27.900 ;
        RECT 138.600 27.200 139.000 27.400 ;
        RECT 140.600 27.200 140.900 27.900 ;
        RECT 135.100 26.900 136.000 27.100 ;
        RECT 138.200 26.900 139.000 27.200 ;
        RECT 135.100 26.800 135.900 26.900 ;
        RECT 138.200 26.800 138.600 26.900 ;
        RECT 139.700 26.800 141.000 27.200 ;
        RECT 131.000 26.600 131.300 26.800 ;
        RECT 130.900 26.200 131.300 26.600 ;
        RECT 127.800 25.400 128.200 26.200 ;
        RECT 128.600 26.100 129.000 26.200 ;
        RECT 128.600 25.800 129.400 26.100 ;
        RECT 130.200 25.800 130.600 26.200 ;
        RECT 129.000 25.600 129.400 25.800 ;
        RECT 130.300 25.700 130.600 25.800 ;
        RECT 130.300 25.400 131.300 25.700 ;
        RECT 131.800 25.400 132.200 26.200 ;
        RECT 132.600 25.400 133.000 26.200 ;
        RECT 133.400 26.100 133.700 26.800 ;
        RECT 134.200 26.100 134.600 26.200 ;
        RECT 133.400 25.800 134.600 26.100 ;
        RECT 131.000 25.200 131.300 25.400 ;
        RECT 117.400 24.800 117.800 24.900 ;
        RECT 115.500 22.200 115.900 24.800 ;
        RECT 117.500 24.500 117.800 24.800 ;
        RECT 124.300 24.800 124.800 25.100 ;
        RECT 125.100 24.800 125.800 25.100 ;
        RECT 118.300 24.500 120.100 24.600 ;
        RECT 115.500 21.800 116.200 22.200 ;
        RECT 115.500 21.100 115.900 21.800 ;
        RECT 116.600 21.500 117.000 24.500 ;
        RECT 117.400 21.700 117.800 24.500 ;
        RECT 118.200 24.300 120.100 24.500 ;
        RECT 116.700 21.400 117.000 21.500 ;
        RECT 118.200 21.500 118.600 24.300 ;
        RECT 119.800 24.100 120.100 24.300 ;
        RECT 120.700 24.400 122.500 24.700 ;
        RECT 120.700 24.100 121.000 24.400 ;
        RECT 118.200 21.400 118.500 21.500 ;
        RECT 116.700 21.100 118.500 21.400 ;
        RECT 119.000 21.400 119.400 24.000 ;
        RECT 119.800 21.700 120.200 24.100 ;
        RECT 120.600 21.400 121.000 24.100 ;
        RECT 119.000 21.100 121.000 21.400 ;
        RECT 122.200 24.100 122.500 24.400 ;
        RECT 122.200 21.100 122.600 24.100 ;
        RECT 124.300 21.100 124.700 24.800 ;
        RECT 125.100 24.200 125.400 24.800 ;
        RECT 127.000 24.700 127.900 25.100 ;
        RECT 125.000 23.800 125.400 24.200 ;
        RECT 127.500 21.100 127.900 24.700 ;
        RECT 128.600 24.800 130.600 25.100 ;
        RECT 128.600 21.100 129.000 24.800 ;
        RECT 130.200 21.400 130.600 24.800 ;
        RECT 131.000 21.700 131.400 25.200 ;
        RECT 133.400 25.100 133.700 25.800 ;
        RECT 135.100 25.200 135.400 26.800 ;
        RECT 136.200 25.800 137.000 26.200 ;
        RECT 139.000 25.800 139.400 26.600 ;
        RECT 139.700 26.200 140.000 26.800 ;
        RECT 139.700 25.800 140.200 26.200 ;
        RECT 131.800 21.400 132.200 25.100 ;
        RECT 130.200 21.100 132.200 21.400 ;
        RECT 132.900 24.700 133.800 25.100 ;
        RECT 135.000 24.800 135.400 25.200 ;
        RECT 137.400 24.800 137.800 25.600 ;
        RECT 139.700 25.100 140.000 25.800 ;
        RECT 140.600 25.100 141.000 25.200 ;
        RECT 139.500 24.800 140.000 25.100 ;
        RECT 140.300 24.800 141.000 25.100 ;
        RECT 132.900 21.100 133.300 24.700 ;
        RECT 135.100 23.500 135.400 24.800 ;
        RECT 135.800 23.800 136.200 24.600 ;
        RECT 136.600 23.800 137.000 24.200 ;
        RECT 136.600 23.500 136.900 23.800 ;
        RECT 135.100 23.200 136.900 23.500 ;
        RECT 135.100 23.100 135.400 23.200 ;
        RECT 135.000 21.100 135.400 23.100 ;
        RECT 136.600 23.100 136.900 23.200 ;
        RECT 136.600 21.100 137.000 23.100 ;
        RECT 139.500 21.100 139.900 24.800 ;
        RECT 140.300 24.200 140.600 24.800 ;
        RECT 141.400 24.400 141.800 25.200 ;
        RECT 140.200 23.800 140.600 24.200 ;
        RECT 142.200 21.100 142.600 27.900 ;
        RECT 143.000 26.800 143.400 27.600 ;
        RECT 145.600 27.100 146.000 29.900 ;
        RECT 147.000 27.900 147.400 29.900 ;
        RECT 147.800 28.000 148.200 29.900 ;
        RECT 149.400 28.000 149.800 29.900 ;
        RECT 147.800 27.900 149.800 28.000 ;
        RECT 147.100 27.200 147.400 27.900 ;
        RECT 147.900 27.700 149.700 27.900 ;
        RECT 149.000 27.200 149.400 27.400 ;
        RECT 145.600 26.900 146.500 27.100 ;
        RECT 145.700 26.800 146.500 26.900 ;
        RECT 147.000 26.800 148.300 27.200 ;
        RECT 149.000 26.900 149.800 27.200 ;
        RECT 149.400 26.800 149.800 26.900 ;
        RECT 144.600 25.800 145.400 26.200 ;
        RECT 143.800 24.800 144.200 25.600 ;
        RECT 146.200 25.200 146.500 26.800 ;
        RECT 146.200 24.800 146.600 25.200 ;
        RECT 147.000 25.100 147.400 25.200 ;
        RECT 148.000 25.100 148.300 26.800 ;
        RECT 148.600 25.800 149.000 26.600 ;
        RECT 147.000 24.800 147.700 25.100 ;
        RECT 148.000 24.800 148.500 25.100 ;
        RECT 145.400 23.800 145.800 24.600 ;
        RECT 146.200 23.500 146.500 24.800 ;
        RECT 147.400 24.200 147.700 24.800 ;
        RECT 147.400 23.800 147.800 24.200 ;
        RECT 144.700 23.200 146.500 23.500 ;
        RECT 144.600 21.100 145.000 23.200 ;
        RECT 146.200 23.100 146.500 23.200 ;
        RECT 146.200 21.100 146.600 23.100 ;
        RECT 148.100 21.100 148.500 24.800 ;
        RECT 0.600 15.700 1.000 19.900 ;
        RECT 2.800 18.200 3.200 19.900 ;
        RECT 2.200 17.900 3.200 18.200 ;
        RECT 5.000 17.900 5.400 19.900 ;
        RECT 7.100 17.900 7.700 19.900 ;
        RECT 2.200 17.500 2.600 17.900 ;
        RECT 5.000 17.600 5.300 17.900 ;
        RECT 3.900 17.300 5.700 17.600 ;
        RECT 7.000 17.500 7.400 17.900 ;
        RECT 3.900 17.200 4.300 17.300 ;
        RECT 5.300 17.200 5.700 17.300 ;
        RECT 2.200 16.500 2.600 16.600 ;
        RECT 4.500 16.500 4.900 16.600 ;
        RECT 2.200 16.200 4.900 16.500 ;
        RECT 5.200 16.500 6.300 16.800 ;
        RECT 5.200 15.900 5.500 16.500 ;
        RECT 5.900 16.400 6.300 16.500 ;
        RECT 7.100 16.600 7.800 17.000 ;
        RECT 7.100 16.100 7.400 16.600 ;
        RECT 3.100 15.700 5.500 15.900 ;
        RECT 0.600 15.600 5.500 15.700 ;
        RECT 6.200 15.800 7.400 16.100 ;
        RECT 0.600 15.500 3.500 15.600 ;
        RECT 0.600 15.400 3.400 15.500 ;
        RECT 6.200 15.200 6.500 15.800 ;
        RECT 9.400 15.600 9.800 19.900 ;
        RECT 7.700 15.300 9.800 15.600 ;
        RECT 7.700 15.200 8.100 15.300 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 8.500 14.900 8.900 15.000 ;
        RECT 2.500 14.200 2.900 14.300 ;
        RECT 6.200 14.200 6.500 14.800 ;
        RECT 7.000 14.600 8.900 14.900 ;
        RECT 7.000 14.500 7.400 14.600 ;
        RECT 1.000 13.900 6.500 14.200 ;
        RECT 1.000 13.800 1.800 13.900 ;
        RECT 0.600 11.100 1.000 13.500 ;
        RECT 3.100 12.800 3.400 13.900 ;
        RECT 5.900 13.800 6.300 13.900 ;
        RECT 9.400 13.600 9.800 15.300 ;
        RECT 7.900 13.300 9.800 13.600 ;
        RECT 7.900 13.200 8.300 13.300 ;
        RECT 2.200 12.100 2.600 12.500 ;
        RECT 3.000 12.400 3.400 12.800 ;
        RECT 3.900 12.700 4.300 12.800 ;
        RECT 3.900 12.400 5.300 12.700 ;
        RECT 5.000 12.100 5.300 12.400 ;
        RECT 7.000 12.100 7.400 12.500 ;
        RECT 2.200 11.800 3.200 12.100 ;
        RECT 2.800 11.100 3.200 11.800 ;
        RECT 5.000 11.100 5.400 12.100 ;
        RECT 7.000 11.800 7.700 12.100 ;
        RECT 7.100 11.100 7.700 11.800 ;
        RECT 9.400 11.100 9.800 13.300 ;
        RECT 11.000 11.100 11.400 19.900 ;
        RECT 11.800 16.200 12.200 19.900 ;
        RECT 12.500 16.200 12.900 16.300 ;
        RECT 11.800 15.900 12.900 16.200 ;
        RECT 14.000 16.200 14.800 19.900 ;
        RECT 15.800 16.200 16.200 16.300 ;
        RECT 16.600 16.200 17.000 19.900 ;
        RECT 14.000 15.900 15.000 16.200 ;
        RECT 15.800 15.900 17.000 16.200 ;
        RECT 12.600 15.600 12.900 15.900 ;
        RECT 12.600 15.300 14.300 15.600 ;
        RECT 13.900 15.200 14.300 15.300 ;
        RECT 14.700 15.200 15.000 15.900 ;
        RECT 17.400 15.700 17.800 19.900 ;
        RECT 19.600 18.200 20.000 19.900 ;
        RECT 19.000 17.900 20.000 18.200 ;
        RECT 21.800 17.900 22.200 19.900 ;
        RECT 23.900 17.900 24.500 19.900 ;
        RECT 19.000 17.500 19.400 17.900 ;
        RECT 21.800 17.600 22.100 17.900 ;
        RECT 20.700 17.300 22.500 17.600 ;
        RECT 23.800 17.500 24.200 17.900 ;
        RECT 20.700 17.200 21.100 17.300 ;
        RECT 22.100 17.200 22.500 17.300 ;
        RECT 19.000 16.500 19.400 16.600 ;
        RECT 21.300 16.500 21.700 16.600 ;
        RECT 19.000 16.200 21.700 16.500 ;
        RECT 22.000 16.500 23.100 16.800 ;
        RECT 22.000 15.900 22.300 16.500 ;
        RECT 22.700 16.400 23.100 16.500 ;
        RECT 23.900 16.600 24.600 17.000 ;
        RECT 23.900 16.100 24.200 16.600 ;
        RECT 19.900 15.700 22.300 15.900 ;
        RECT 17.400 15.600 22.300 15.700 ;
        RECT 23.000 15.800 24.200 16.100 ;
        RECT 17.400 15.500 20.300 15.600 ;
        RECT 17.400 15.400 20.200 15.500 ;
        RECT 12.800 14.900 13.200 15.000 ;
        RECT 14.700 14.900 15.400 15.200 ;
        RECT 12.800 14.600 14.100 14.900 ;
        RECT 13.800 14.300 14.100 14.600 ;
        RECT 14.500 14.800 15.400 14.900 ;
        RECT 14.500 14.600 15.000 14.800 ;
        RECT 13.800 13.900 14.200 14.300 ;
        RECT 12.500 13.400 12.900 13.500 ;
        RECT 11.800 13.100 12.900 13.400 ;
        RECT 11.800 11.100 12.200 13.100 ;
        RECT 14.500 12.900 14.800 14.600 ;
        RECT 19.300 14.200 19.700 14.300 ;
        RECT 23.000 14.200 23.300 15.800 ;
        RECT 26.200 15.600 26.600 19.900 ;
        RECT 27.000 16.200 27.400 19.900 ;
        RECT 29.200 19.200 30.000 19.900 ;
        RECT 29.200 18.800 30.600 19.200 ;
        RECT 27.700 16.200 28.100 16.300 ;
        RECT 27.000 15.900 28.100 16.200 ;
        RECT 29.200 16.200 30.000 18.800 ;
        RECT 31.000 16.200 31.400 16.300 ;
        RECT 31.800 16.200 32.200 19.900 ;
        RECT 29.200 15.900 30.200 16.200 ;
        RECT 31.000 15.900 32.200 16.200 ;
        RECT 24.500 15.300 26.600 15.600 ;
        RECT 27.800 15.600 28.100 15.900 ;
        RECT 27.800 15.300 29.500 15.600 ;
        RECT 24.500 15.200 24.900 15.300 ;
        RECT 25.300 14.900 25.700 15.000 ;
        RECT 23.800 14.600 25.700 14.900 ;
        RECT 23.800 14.500 24.200 14.600 ;
        RECT 17.800 13.900 23.300 14.200 ;
        RECT 17.800 13.800 18.600 13.900 ;
        RECT 15.800 13.400 16.200 13.500 ;
        RECT 15.800 13.100 17.000 13.400 ;
        RECT 14.000 12.200 14.800 12.900 ;
        RECT 13.400 11.800 14.800 12.200 ;
        RECT 14.000 11.100 14.800 11.800 ;
        RECT 16.600 11.100 17.000 13.100 ;
        RECT 17.400 11.100 17.800 13.500 ;
        RECT 19.900 12.800 20.200 13.900 ;
        RECT 20.600 13.800 21.000 13.900 ;
        RECT 22.700 13.800 23.100 13.900 ;
        RECT 26.200 13.600 26.600 15.300 ;
        RECT 29.100 15.200 29.500 15.300 ;
        RECT 29.900 15.200 30.200 15.900 ;
        RECT 32.600 15.700 33.000 19.900 ;
        RECT 34.800 18.200 35.200 19.900 ;
        RECT 34.200 17.900 35.200 18.200 ;
        RECT 37.000 17.900 37.400 19.900 ;
        RECT 39.100 17.900 39.700 19.900 ;
        RECT 34.200 17.500 34.600 17.900 ;
        RECT 37.000 17.600 37.300 17.900 ;
        RECT 35.900 17.300 37.700 17.600 ;
        RECT 39.000 17.500 39.400 17.900 ;
        RECT 35.900 17.200 36.300 17.300 ;
        RECT 37.300 17.200 37.700 17.300 ;
        RECT 34.200 16.500 34.600 16.600 ;
        RECT 36.500 16.500 36.900 16.600 ;
        RECT 34.200 16.200 36.900 16.500 ;
        RECT 37.200 16.500 38.300 16.800 ;
        RECT 37.200 15.900 37.500 16.500 ;
        RECT 37.900 16.400 38.300 16.500 ;
        RECT 39.100 16.600 39.800 17.000 ;
        RECT 39.100 16.100 39.400 16.600 ;
        RECT 35.100 15.700 37.500 15.900 ;
        RECT 32.600 15.600 37.500 15.700 ;
        RECT 38.200 15.800 39.400 16.100 ;
        RECT 32.600 15.500 35.500 15.600 ;
        RECT 32.600 15.400 35.400 15.500 ;
        RECT 28.000 14.900 28.400 15.000 ;
        RECT 29.900 14.900 30.600 15.200 ;
        RECT 35.800 15.100 36.200 15.200 ;
        RECT 36.600 15.100 37.000 15.200 ;
        RECT 28.000 14.600 29.300 14.900 ;
        RECT 29.000 14.300 29.300 14.600 ;
        RECT 29.700 14.800 30.600 14.900 ;
        RECT 33.700 14.800 37.000 15.100 ;
        RECT 29.700 14.600 30.200 14.800 ;
        RECT 33.700 14.700 34.100 14.800 ;
        RECT 27.000 14.100 27.800 14.200 ;
        RECT 27.000 13.800 28.700 14.100 ;
        RECT 29.000 13.900 29.400 14.300 ;
        RECT 24.700 13.300 26.600 13.600 ;
        RECT 28.400 13.600 28.700 13.800 ;
        RECT 27.700 13.400 28.100 13.500 ;
        RECT 24.700 13.200 25.100 13.300 ;
        RECT 19.000 12.100 19.400 12.500 ;
        RECT 19.800 12.400 20.200 12.800 ;
        RECT 20.700 12.700 21.100 12.800 ;
        RECT 20.700 12.400 22.100 12.700 ;
        RECT 21.800 12.100 22.100 12.400 ;
        RECT 23.800 12.100 24.200 12.500 ;
        RECT 19.000 11.800 20.000 12.100 ;
        RECT 19.600 11.100 20.000 11.800 ;
        RECT 21.800 11.100 22.200 12.100 ;
        RECT 23.800 11.800 24.500 12.100 ;
        RECT 23.900 11.100 24.500 11.800 ;
        RECT 26.200 11.100 26.600 13.300 ;
        RECT 27.000 13.100 28.100 13.400 ;
        RECT 28.400 13.300 29.400 13.600 ;
        RECT 28.600 13.200 29.400 13.300 ;
        RECT 27.000 11.100 27.400 13.100 ;
        RECT 29.700 12.900 30.000 14.600 ;
        RECT 34.500 14.200 34.900 14.300 ;
        RECT 38.200 14.200 38.500 15.800 ;
        RECT 41.400 15.600 41.800 19.900 ;
        RECT 39.700 15.300 41.800 15.600 ;
        RECT 39.700 15.200 40.100 15.300 ;
        RECT 40.500 14.900 40.900 15.000 ;
        RECT 39.000 14.600 40.900 14.900 ;
        RECT 39.000 14.500 39.400 14.600 ;
        RECT 30.400 13.800 30.800 14.200 ;
        RECT 31.400 13.800 32.200 14.200 ;
        RECT 33.000 13.900 38.500 14.200 ;
        RECT 33.000 13.800 33.800 13.900 ;
        RECT 30.400 13.600 30.700 13.800 ;
        RECT 30.300 13.200 30.700 13.600 ;
        RECT 31.000 13.400 31.400 13.500 ;
        RECT 31.000 13.100 32.200 13.400 ;
        RECT 29.200 11.100 30.000 12.900 ;
        RECT 31.800 11.100 32.200 13.100 ;
        RECT 32.600 11.100 33.000 13.500 ;
        RECT 35.100 12.800 35.400 13.900 ;
        RECT 37.900 13.800 38.300 13.900 ;
        RECT 41.400 13.600 41.800 15.300 ;
        RECT 39.900 13.300 41.800 13.600 ;
        RECT 39.900 13.200 40.300 13.300 ;
        RECT 34.200 12.100 34.600 12.500 ;
        RECT 35.000 12.400 35.400 12.800 ;
        RECT 35.900 12.700 36.300 12.800 ;
        RECT 35.900 12.400 37.300 12.700 ;
        RECT 37.000 12.100 37.300 12.400 ;
        RECT 39.000 12.100 39.400 12.500 ;
        RECT 34.200 11.800 35.200 12.100 ;
        RECT 34.800 11.100 35.200 11.800 ;
        RECT 37.000 11.100 37.400 12.100 ;
        RECT 39.000 11.800 39.700 12.100 ;
        RECT 39.100 11.100 39.700 11.800 ;
        RECT 41.400 11.100 41.800 13.300 ;
        RECT 42.200 15.800 42.600 19.900 ;
        RECT 43.800 17.900 44.200 19.900 ;
        RECT 43.800 15.800 44.100 17.900 ;
        RECT 45.700 16.300 46.100 19.900 ;
        RECT 49.100 16.300 49.500 19.900 ;
        RECT 45.700 15.900 46.600 16.300 ;
        RECT 48.600 15.900 49.500 16.300 ;
        RECT 42.200 15.200 42.500 15.800 ;
        RECT 42.900 15.500 44.100 15.800 ;
        RECT 42.200 14.800 42.600 15.200 ;
        RECT 42.200 13.100 42.500 14.800 ;
        RECT 42.900 13.800 43.200 15.500 ;
        RECT 43.800 14.800 44.200 15.200 ;
        RECT 45.400 14.800 45.800 15.600 ;
        RECT 43.800 14.400 44.100 14.800 ;
        RECT 43.600 14.100 44.100 14.400 ;
        RECT 44.600 14.100 45.000 14.600 ;
        RECT 46.200 14.200 46.500 15.900 ;
        RECT 47.800 15.100 48.200 15.200 ;
        RECT 48.700 15.100 49.000 15.900 ;
        RECT 51.800 15.700 52.200 19.900 ;
        RECT 54.000 18.200 54.400 19.900 ;
        RECT 53.400 17.900 54.400 18.200 ;
        RECT 56.200 17.900 56.600 19.900 ;
        RECT 58.300 17.900 58.900 19.900 ;
        RECT 53.400 17.500 53.800 17.900 ;
        RECT 56.200 17.600 56.500 17.900 ;
        RECT 55.100 17.300 56.900 17.600 ;
        RECT 58.200 17.500 58.600 17.900 ;
        RECT 55.100 17.200 55.500 17.300 ;
        RECT 56.500 17.200 56.900 17.300 ;
        RECT 53.400 16.500 53.800 16.600 ;
        RECT 55.700 16.500 56.100 16.600 ;
        RECT 53.400 16.200 56.100 16.500 ;
        RECT 56.400 16.500 57.500 16.800 ;
        RECT 56.400 15.900 56.700 16.500 ;
        RECT 57.100 16.400 57.500 16.500 ;
        RECT 58.300 16.600 59.000 17.000 ;
        RECT 58.300 16.100 58.600 16.600 ;
        RECT 54.300 15.700 56.700 15.900 ;
        RECT 51.800 15.600 56.700 15.700 ;
        RECT 57.400 15.800 58.600 16.100 ;
        RECT 47.800 14.800 49.000 15.100 ;
        RECT 49.400 14.800 49.800 15.600 ;
        RECT 51.800 15.500 54.700 15.600 ;
        RECT 51.800 15.400 54.600 15.500 ;
        RECT 57.400 15.200 57.700 15.800 ;
        RECT 60.600 15.600 61.000 19.900 ;
        RECT 58.900 15.300 61.000 15.600 ;
        RECT 61.400 15.700 61.800 19.900 ;
        RECT 63.600 18.200 64.000 19.900 ;
        RECT 63.000 17.900 64.000 18.200 ;
        RECT 65.800 17.900 66.200 19.900 ;
        RECT 67.900 17.900 68.500 19.900 ;
        RECT 63.000 17.500 63.400 17.900 ;
        RECT 65.800 17.600 66.100 17.900 ;
        RECT 64.700 17.300 66.500 17.600 ;
        RECT 67.800 17.500 68.200 17.900 ;
        RECT 64.700 17.200 65.100 17.300 ;
        RECT 66.100 17.200 66.500 17.300 ;
        RECT 63.000 16.500 63.400 16.600 ;
        RECT 65.300 16.500 65.700 16.600 ;
        RECT 63.000 16.200 65.700 16.500 ;
        RECT 66.000 16.500 67.100 16.800 ;
        RECT 66.000 15.900 66.300 16.500 ;
        RECT 66.700 16.400 67.100 16.500 ;
        RECT 67.900 16.600 68.600 17.000 ;
        RECT 67.900 16.100 68.200 16.600 ;
        RECT 63.900 15.700 66.300 15.900 ;
        RECT 61.400 15.600 66.300 15.700 ;
        RECT 67.000 15.800 68.200 16.100 ;
        RECT 61.400 15.500 64.300 15.600 ;
        RECT 61.400 15.400 64.200 15.500 ;
        RECT 58.900 15.200 59.300 15.300 ;
        RECT 55.000 15.100 55.400 15.200 ;
        RECT 52.900 14.800 55.400 15.100 ;
        RECT 57.400 14.800 57.800 15.200 ;
        RECT 59.700 14.900 60.100 15.000 ;
        RECT 48.700 14.200 49.000 14.800 ;
        RECT 52.900 14.700 53.300 14.800 ;
        RECT 54.200 14.700 54.600 14.800 ;
        RECT 53.700 14.200 54.100 14.300 ;
        RECT 57.400 14.200 57.700 14.800 ;
        RECT 58.200 14.600 60.100 14.900 ;
        RECT 58.200 14.500 58.600 14.600 ;
        RECT 45.400 14.100 45.800 14.200 ;
        RECT 43.600 14.000 44.000 14.100 ;
        RECT 44.600 13.800 45.800 14.100 ;
        RECT 46.200 14.100 46.600 14.200 ;
        RECT 46.200 13.800 48.100 14.100 ;
        RECT 48.600 13.800 49.000 14.200 ;
        RECT 52.200 13.900 57.700 14.200 ;
        RECT 52.200 13.800 53.000 13.900 ;
        RECT 42.800 13.700 43.200 13.800 ;
        RECT 42.800 13.500 44.300 13.700 ;
        RECT 42.800 13.400 44.900 13.500 ;
        RECT 44.000 13.200 44.900 13.400 ;
        RECT 44.600 13.100 44.900 13.200 ;
        RECT 42.200 12.600 42.900 13.100 ;
        RECT 42.500 11.100 42.900 12.600 ;
        RECT 44.600 11.100 45.000 13.100 ;
        RECT 46.200 12.100 46.500 13.800 ;
        RECT 47.800 13.200 48.100 13.800 ;
        RECT 47.000 12.400 47.400 13.200 ;
        RECT 47.800 12.400 48.200 13.200 ;
        RECT 48.700 12.100 49.000 13.800 ;
        RECT 46.200 11.100 46.600 12.100 ;
        RECT 48.600 11.100 49.000 12.100 ;
        RECT 51.800 11.100 52.200 13.500 ;
        RECT 54.300 13.200 54.600 13.900 ;
        RECT 57.100 13.800 57.500 13.900 ;
        RECT 60.600 13.600 61.000 15.300 ;
        RECT 64.600 15.100 65.000 15.200 ;
        RECT 62.500 14.800 65.000 15.100 ;
        RECT 62.500 14.700 62.900 14.800 ;
        RECT 63.300 14.200 63.700 14.300 ;
        RECT 67.000 14.200 67.300 15.800 ;
        RECT 70.200 15.600 70.600 19.900 ;
        RECT 68.500 15.300 70.600 15.600 ;
        RECT 68.500 15.200 68.900 15.300 ;
        RECT 69.300 14.900 69.700 15.000 ;
        RECT 67.800 14.600 69.700 14.900 ;
        RECT 67.800 14.500 68.200 14.600 ;
        RECT 61.800 13.900 67.300 14.200 ;
        RECT 61.800 13.800 62.600 13.900 ;
        RECT 63.800 13.800 64.200 13.900 ;
        RECT 66.700 13.800 67.100 13.900 ;
        RECT 59.100 13.300 61.000 13.600 ;
        RECT 59.100 13.200 59.500 13.300 ;
        RECT 53.400 12.100 53.800 12.500 ;
        RECT 54.200 12.400 54.600 13.200 ;
        RECT 55.100 12.700 55.500 12.800 ;
        RECT 55.100 12.400 56.500 12.700 ;
        RECT 56.200 12.100 56.500 12.400 ;
        RECT 58.200 12.100 58.600 12.500 ;
        RECT 53.400 11.800 54.400 12.100 ;
        RECT 54.000 11.100 54.400 11.800 ;
        RECT 56.200 11.100 56.600 12.100 ;
        RECT 58.200 11.800 58.900 12.100 ;
        RECT 58.300 11.100 58.900 11.800 ;
        RECT 60.600 11.100 61.000 13.300 ;
        RECT 61.400 11.100 61.800 13.500 ;
        RECT 63.900 12.800 64.200 13.800 ;
        RECT 70.200 13.600 70.600 15.300 ;
        RECT 71.800 15.100 72.200 19.900 ;
        RECT 72.600 15.800 73.000 17.200 ;
        RECT 73.700 16.300 74.100 19.900 ;
        RECT 73.700 15.900 74.600 16.300 ;
        RECT 73.400 15.100 73.800 15.600 ;
        RECT 71.800 14.800 73.800 15.100 ;
        RECT 68.700 13.300 70.600 13.600 ;
        RECT 71.000 13.400 71.400 14.200 ;
        RECT 68.700 13.200 69.100 13.300 ;
        RECT 63.000 12.100 63.400 12.500 ;
        RECT 63.800 12.400 64.200 12.800 ;
        RECT 64.700 12.700 65.100 12.800 ;
        RECT 64.700 12.400 66.100 12.700 ;
        RECT 65.800 12.100 66.100 12.400 ;
        RECT 67.800 12.100 68.200 12.500 ;
        RECT 63.000 11.800 64.000 12.100 ;
        RECT 63.600 11.100 64.000 11.800 ;
        RECT 65.800 11.100 66.200 12.100 ;
        RECT 67.800 11.800 68.500 12.100 ;
        RECT 67.900 11.100 68.500 11.800 ;
        RECT 70.200 11.100 70.600 13.300 ;
        RECT 71.800 13.100 72.200 14.800 ;
        RECT 73.400 14.200 73.700 14.800 ;
        RECT 74.200 14.200 74.500 15.900 ;
        RECT 73.400 13.800 73.800 14.200 ;
        RECT 74.200 14.100 74.600 14.200 ;
        RECT 74.200 13.800 76.100 14.100 ;
        RECT 71.800 12.800 72.700 13.100 ;
        RECT 72.300 11.100 72.700 12.800 ;
        RECT 74.200 12.100 74.500 13.800 ;
        RECT 75.800 13.200 76.100 13.800 ;
        RECT 75.000 12.400 75.400 13.200 ;
        RECT 75.800 12.400 76.200 13.200 ;
        RECT 74.200 11.100 74.600 12.100 ;
        RECT 76.600 11.100 77.000 19.900 ;
        RECT 78.700 16.200 79.100 19.900 ;
        RECT 79.400 16.800 79.800 17.200 ;
        RECT 79.500 16.200 79.800 16.800 ;
        RECT 80.900 16.300 81.300 19.900 ;
        RECT 78.700 15.900 79.200 16.200 ;
        RECT 79.500 15.900 80.200 16.200 ;
        RECT 80.900 15.900 81.800 16.300 ;
        RECT 83.000 15.900 83.400 19.900 ;
        RECT 84.600 17.900 85.000 19.900 ;
        RECT 78.200 14.400 78.600 15.200 ;
        RECT 78.900 14.200 79.200 15.900 ;
        RECT 79.800 15.800 80.200 15.900 ;
        RECT 79.800 15.100 80.100 15.800 ;
        RECT 80.600 15.100 81.000 15.600 ;
        RECT 79.800 14.800 81.000 15.100 ;
        RECT 81.400 14.200 81.700 15.900 ;
        RECT 83.000 15.200 83.300 15.900 ;
        RECT 84.600 15.800 84.900 17.900 ;
        RECT 83.700 15.500 84.900 15.800 ;
        RECT 86.200 15.900 86.600 19.900 ;
        RECT 87.800 17.900 88.200 19.900 ;
        RECT 82.200 14.800 82.600 15.200 ;
        RECT 83.000 14.800 83.400 15.200 ;
        RECT 77.400 14.100 77.800 14.200 ;
        RECT 77.400 13.800 78.200 14.100 ;
        RECT 78.900 13.800 80.200 14.200 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 82.200 14.100 82.500 14.800 ;
        RECT 81.400 13.800 82.500 14.100 ;
        RECT 77.800 13.600 78.200 13.800 ;
        RECT 77.500 13.100 79.300 13.300 ;
        RECT 79.800 13.100 80.100 13.800 ;
        RECT 77.400 13.000 79.400 13.100 ;
        RECT 77.400 11.100 77.800 13.000 ;
        RECT 79.000 11.100 79.400 13.000 ;
        RECT 79.800 11.100 80.200 13.100 ;
        RECT 81.400 12.100 81.700 13.800 ;
        RECT 82.200 12.400 82.600 13.200 ;
        RECT 83.000 13.100 83.300 14.800 ;
        RECT 83.700 13.800 84.000 15.500 ;
        RECT 86.200 15.200 86.500 15.900 ;
        RECT 87.800 15.800 88.100 17.900 ;
        RECT 86.900 15.500 88.100 15.800 ;
        RECT 84.600 14.800 85.000 15.200 ;
        RECT 86.200 14.800 86.600 15.200 ;
        RECT 84.600 14.400 84.900 14.800 ;
        RECT 84.400 14.100 84.900 14.400 ;
        RECT 84.400 14.000 84.800 14.100 ;
        RECT 85.400 13.800 85.800 14.600 ;
        RECT 83.600 13.700 84.000 13.800 ;
        RECT 83.600 13.500 85.100 13.700 ;
        RECT 83.600 13.400 85.700 13.500 ;
        RECT 84.800 13.200 85.700 13.400 ;
        RECT 85.400 13.100 85.700 13.200 ;
        RECT 86.200 13.100 86.500 14.800 ;
        RECT 86.900 13.800 87.200 15.500 ;
        RECT 87.800 14.800 88.200 15.200 ;
        RECT 87.800 14.400 88.100 14.800 ;
        RECT 87.600 14.000 88.200 14.400 ;
        RECT 88.600 14.100 89.000 14.600 ;
        RECT 89.400 14.100 89.800 19.900 ;
        RECT 91.000 15.900 91.400 19.900 ;
        RECT 91.800 16.200 92.200 19.900 ;
        RECT 93.400 16.200 93.800 19.900 ;
        RECT 95.000 17.900 95.400 19.900 ;
        RECT 95.100 17.800 95.400 17.900 ;
        RECT 96.600 17.900 97.000 19.900 ;
        RECT 96.600 17.800 96.900 17.900 ;
        RECT 95.100 17.500 96.900 17.800 ;
        RECT 95.800 16.400 96.200 17.200 ;
        RECT 96.600 16.200 96.900 17.500 ;
        RECT 98.700 16.300 99.100 19.900 ;
        RECT 91.800 15.900 93.800 16.200 ;
        RECT 91.100 15.200 91.400 15.900 ;
        RECT 94.200 15.400 94.600 16.200 ;
        RECT 96.600 15.800 97.000 16.200 ;
        RECT 98.200 15.900 99.100 16.300 ;
        RECT 101.400 17.100 101.800 19.900 ;
        RECT 103.000 17.900 103.400 19.900 ;
        RECT 103.100 17.800 103.400 17.900 ;
        RECT 104.600 17.900 105.000 19.900 ;
        RECT 104.600 17.800 104.900 17.900 ;
        RECT 103.100 17.500 104.900 17.800 ;
        RECT 101.400 16.800 102.500 17.100 ;
        RECT 93.000 15.200 93.400 15.400 ;
        RECT 91.000 14.900 92.200 15.200 ;
        RECT 93.000 14.900 93.800 15.200 ;
        RECT 91.000 14.800 91.400 14.900 ;
        RECT 88.600 13.800 89.800 14.100 ;
        RECT 86.800 13.700 87.200 13.800 ;
        RECT 86.800 13.500 88.300 13.700 ;
        RECT 86.800 13.400 88.900 13.500 ;
        RECT 88.000 13.200 88.900 13.400 ;
        RECT 88.600 13.100 88.900 13.200 ;
        RECT 83.000 12.600 83.700 13.100 ;
        RECT 83.300 12.200 83.700 12.600 ;
        RECT 81.400 11.100 81.800 12.100 ;
        RECT 83.000 11.800 83.700 12.200 ;
        RECT 83.300 11.100 83.700 11.800 ;
        RECT 85.400 11.100 85.800 13.100 ;
        RECT 86.200 12.600 86.900 13.100 ;
        RECT 86.500 12.200 86.900 12.600 ;
        RECT 86.200 11.800 86.900 12.200 ;
        RECT 86.500 11.100 86.900 11.800 ;
        RECT 88.600 11.100 89.000 13.100 ;
        RECT 89.400 11.100 89.800 13.800 ;
        RECT 91.900 13.200 92.200 14.900 ;
        RECT 93.400 14.800 93.800 14.900 ;
        RECT 95.000 14.800 95.800 15.200 ;
        RECT 92.600 13.800 93.000 14.600 ;
        RECT 96.600 14.200 96.900 15.800 ;
        RECT 96.100 14.100 96.900 14.200 ;
        RECT 97.400 14.800 97.800 15.200 ;
        RECT 97.400 14.100 97.700 14.800 ;
        RECT 98.300 14.200 98.600 15.900 ;
        RECT 99.000 15.100 99.400 15.600 ;
        RECT 101.400 15.100 101.800 16.800 ;
        RECT 102.200 16.200 102.500 16.800 ;
        RECT 103.100 16.200 103.400 17.500 ;
        RECT 103.800 16.400 104.200 17.200 ;
        RECT 102.200 15.800 102.600 16.200 ;
        RECT 103.000 15.800 103.400 16.200 ;
        RECT 99.000 14.800 101.800 15.100 ;
        RECT 96.000 13.800 97.700 14.100 ;
        RECT 98.200 13.800 98.600 14.200 ;
        RECT 90.200 13.100 90.600 13.200 ;
        RECT 91.000 13.100 91.400 13.200 ;
        RECT 90.200 12.800 91.400 13.100 ;
        RECT 90.200 12.400 90.600 12.800 ;
        RECT 91.100 12.400 91.500 12.800 ;
        RECT 91.800 11.100 92.200 13.200 ;
        RECT 96.000 11.100 96.400 13.800 ;
        RECT 97.400 12.400 97.800 13.200 ;
        RECT 98.300 12.200 98.600 13.800 ;
        RECT 98.200 11.100 98.600 12.200 ;
        RECT 101.400 11.100 101.800 14.800 ;
        RECT 103.100 14.200 103.400 15.800 ;
        RECT 105.400 15.400 105.800 16.200 ;
        RECT 104.200 14.800 105.000 15.200 ;
        RECT 103.100 14.100 103.900 14.200 ;
        RECT 103.100 13.900 104.000 14.100 ;
        RECT 102.200 12.400 102.600 13.200 ;
        RECT 103.600 11.100 104.000 13.900 ;
        RECT 106.200 11.100 106.600 19.900 ;
        RECT 108.900 17.200 109.300 19.900 ;
        RECT 111.800 17.900 112.200 19.900 ;
        RECT 108.200 16.800 108.600 17.200 ;
        RECT 108.900 16.800 109.800 17.200 ;
        RECT 108.200 16.200 108.500 16.800 ;
        RECT 108.900 16.200 109.300 16.800 ;
        RECT 107.800 15.900 108.500 16.200 ;
        RECT 108.800 15.900 109.300 16.200 ;
        RECT 107.800 15.800 108.200 15.900 ;
        RECT 108.800 14.200 109.100 15.900 ;
        RECT 111.900 15.800 112.200 17.900 ;
        RECT 113.400 15.900 113.800 19.900 ;
        RECT 114.200 16.900 114.600 19.900 ;
        RECT 114.300 16.600 114.600 16.900 ;
        RECT 115.800 19.600 117.800 19.900 ;
        RECT 115.800 16.900 116.200 19.600 ;
        RECT 116.600 16.900 117.000 19.300 ;
        RECT 117.400 17.000 117.800 19.600 ;
        RECT 118.300 19.600 120.100 19.900 ;
        RECT 118.300 19.500 118.600 19.600 ;
        RECT 115.800 16.600 116.100 16.900 ;
        RECT 114.300 16.300 116.100 16.600 ;
        RECT 116.700 16.700 117.000 16.900 ;
        RECT 118.200 16.700 118.600 19.500 ;
        RECT 119.800 19.500 120.100 19.600 ;
        RECT 116.700 16.500 118.600 16.700 ;
        RECT 119.000 16.500 119.400 19.300 ;
        RECT 119.800 16.500 120.200 19.500 ;
        RECT 116.700 16.400 118.500 16.500 ;
        RECT 119.000 16.200 119.300 16.500 ;
        RECT 119.000 16.100 119.400 16.200 ;
        RECT 111.900 15.500 113.100 15.800 ;
        RECT 109.400 14.400 109.800 15.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 107.800 13.800 109.100 14.200 ;
        RECT 110.200 14.100 110.600 14.200 ;
        RECT 109.800 13.800 110.600 14.100 ;
        RECT 111.000 13.800 111.400 14.600 ;
        RECT 111.900 14.400 112.200 14.800 ;
        RECT 111.900 14.100 112.400 14.400 ;
        RECT 112.000 14.000 112.400 14.100 ;
        RECT 112.800 13.800 113.100 15.500 ;
        RECT 113.500 15.200 113.800 15.900 ;
        RECT 117.700 15.800 119.400 16.100 ;
        RECT 120.600 15.900 121.000 19.900 ;
        RECT 121.400 16.200 121.800 19.900 ;
        RECT 123.000 16.200 123.400 19.900 ;
        RECT 125.100 16.300 125.500 19.900 ;
        RECT 127.000 17.900 127.400 19.900 ;
        RECT 127.100 17.800 127.400 17.900 ;
        RECT 128.600 17.900 129.000 19.900 ;
        RECT 128.600 17.800 128.900 17.900 ;
        RECT 127.100 17.500 128.900 17.800 ;
        RECT 126.200 17.100 126.600 17.200 ;
        RECT 127.800 17.100 128.200 17.200 ;
        RECT 126.200 16.800 128.200 17.100 ;
        RECT 127.800 16.400 128.200 16.800 ;
        RECT 121.400 15.900 123.400 16.200 ;
        RECT 124.600 15.900 125.500 16.300 ;
        RECT 128.600 16.200 128.900 17.500 ;
        RECT 129.400 16.200 129.800 19.900 ;
        RECT 131.600 17.200 132.400 19.900 ;
        RECT 131.600 16.800 133.000 17.200 ;
        RECT 130.200 16.200 130.600 16.300 ;
        RECT 131.600 16.200 132.400 16.800 ;
        RECT 113.400 14.800 113.800 15.200 ;
        RECT 116.600 14.800 117.400 15.200 ;
        RECT 107.000 12.400 107.400 13.200 ;
        RECT 107.900 13.100 108.200 13.800 ;
        RECT 109.800 13.600 110.200 13.800 ;
        RECT 112.800 13.700 113.200 13.800 ;
        RECT 111.700 13.500 113.200 13.700 ;
        RECT 111.100 13.400 113.200 13.500 ;
        RECT 108.700 13.100 110.500 13.300 ;
        RECT 111.100 13.200 112.000 13.400 ;
        RECT 111.100 13.100 111.400 13.200 ;
        RECT 113.500 13.100 113.800 14.800 ;
        RECT 115.000 14.100 115.400 14.200 ;
        RECT 115.800 14.100 116.600 14.200 ;
        RECT 115.000 13.800 116.600 14.100 ;
        RECT 107.800 11.100 108.200 13.100 ;
        RECT 108.600 13.000 110.600 13.100 ;
        RECT 108.600 11.100 109.000 13.000 ;
        RECT 110.200 11.100 110.600 13.000 ;
        RECT 111.000 11.100 111.400 13.100 ;
        RECT 113.100 12.600 113.800 13.100 ;
        RECT 114.200 13.100 114.600 13.200 ;
        RECT 115.000 13.100 115.900 13.200 ;
        RECT 114.200 12.800 115.900 13.100 ;
        RECT 117.700 13.100 118.000 15.800 ;
        RECT 120.700 15.200 121.000 15.900 ;
        RECT 122.600 15.200 123.000 15.400 ;
        RECT 120.600 14.900 121.800 15.200 ;
        RECT 122.600 14.900 123.400 15.200 ;
        RECT 120.600 14.800 121.000 14.900 ;
        RECT 121.500 13.200 121.800 14.900 ;
        RECT 123.000 14.800 123.400 14.900 ;
        RECT 122.200 13.800 122.600 14.600 ;
        RECT 124.700 14.200 125.000 15.900 ;
        RECT 125.400 14.800 125.800 15.600 ;
        RECT 126.200 15.400 126.600 16.200 ;
        RECT 128.600 15.800 129.000 16.200 ;
        RECT 129.400 15.900 130.600 16.200 ;
        RECT 131.400 15.900 132.400 16.200 ;
        RECT 133.500 16.200 133.900 16.300 ;
        RECT 134.200 16.200 134.600 19.900 ;
        RECT 133.500 15.900 134.600 16.200 ;
        RECT 127.000 14.800 127.800 15.200 ;
        RECT 128.600 14.200 128.900 15.800 ;
        RECT 131.400 15.200 131.700 15.900 ;
        RECT 133.500 15.600 133.800 15.900 ;
        RECT 132.100 15.300 133.800 15.600 ;
        RECT 135.000 15.700 135.400 19.900 ;
        RECT 137.200 18.200 137.600 19.900 ;
        RECT 136.600 17.900 137.600 18.200 ;
        RECT 139.400 17.900 139.800 19.900 ;
        RECT 141.500 17.900 142.100 19.900 ;
        RECT 136.600 17.500 137.000 17.900 ;
        RECT 139.400 17.600 139.700 17.900 ;
        RECT 138.300 17.300 140.100 17.600 ;
        RECT 141.400 17.500 141.800 17.900 ;
        RECT 138.300 17.200 138.700 17.300 ;
        RECT 139.700 17.200 140.100 17.300 ;
        RECT 136.600 16.500 137.000 16.600 ;
        RECT 138.900 16.500 139.300 16.600 ;
        RECT 136.600 16.200 139.300 16.500 ;
        RECT 139.600 16.500 140.700 16.800 ;
        RECT 139.600 15.900 139.900 16.500 ;
        RECT 140.300 16.400 140.700 16.500 ;
        RECT 141.500 16.600 142.200 17.000 ;
        RECT 141.500 16.100 141.800 16.600 ;
        RECT 137.500 15.700 139.900 15.900 ;
        RECT 135.000 15.600 139.900 15.700 ;
        RECT 140.600 15.800 141.800 16.100 ;
        RECT 135.000 15.500 137.900 15.600 ;
        RECT 135.000 15.400 137.800 15.500 ;
        RECT 132.100 15.200 132.500 15.300 ;
        RECT 131.000 14.900 131.700 15.200 ;
        RECT 138.200 15.100 138.600 15.200 ;
        RECT 133.200 14.900 133.600 15.000 ;
        RECT 131.000 14.800 131.900 14.900 ;
        RECT 131.400 14.600 131.900 14.800 ;
        RECT 124.600 13.800 125.000 14.200 ;
        RECT 128.100 14.100 128.900 14.200 ;
        RECT 129.400 14.100 130.200 14.200 ;
        RECT 120.600 13.100 121.000 13.200 ;
        RECT 117.700 12.800 121.000 13.100 ;
        RECT 113.100 12.200 113.500 12.600 ;
        RECT 117.700 12.500 118.000 12.800 ;
        RECT 116.000 12.200 118.000 12.500 ;
        RECT 120.700 12.400 121.100 12.800 ;
        RECT 113.100 11.800 113.800 12.200 ;
        RECT 116.000 12.100 116.300 12.200 ;
        RECT 115.800 11.800 116.300 12.100 ;
        RECT 117.400 12.100 118.000 12.200 ;
        RECT 113.100 11.100 113.500 11.800 ;
        RECT 115.800 11.100 116.200 11.800 ;
        RECT 117.400 11.100 117.800 12.100 ;
        RECT 121.400 11.100 121.800 13.200 ;
        RECT 123.800 12.400 124.200 13.200 ;
        RECT 124.700 12.200 125.000 13.800 ;
        RECT 124.600 11.100 125.000 12.200 ;
        RECT 128.000 13.800 130.200 14.100 ;
        RECT 130.800 13.800 131.200 14.200 ;
        RECT 128.000 11.100 128.400 13.800 ;
        RECT 130.900 13.600 131.200 13.800 ;
        RECT 130.200 13.400 130.600 13.500 ;
        RECT 129.400 13.100 130.600 13.400 ;
        RECT 130.900 13.200 131.300 13.600 ;
        RECT 129.400 11.100 129.800 13.100 ;
        RECT 131.600 12.900 131.900 14.600 ;
        RECT 132.300 14.600 133.600 14.900 ;
        RECT 136.100 14.800 138.600 15.100 ;
        RECT 136.100 14.700 136.500 14.800 ;
        RECT 137.400 14.700 137.800 14.800 ;
        RECT 132.300 14.300 132.600 14.600 ;
        RECT 132.200 13.900 132.600 14.300 ;
        RECT 136.900 14.200 137.300 14.300 ;
        RECT 140.600 14.200 140.900 15.800 ;
        RECT 143.800 15.600 144.200 19.900 ;
        RECT 144.600 16.200 145.000 19.900 ;
        RECT 148.300 19.200 148.700 19.900 ;
        RECT 147.800 18.800 148.700 19.200 ;
        RECT 148.300 16.200 148.700 18.800 ;
        RECT 149.000 16.800 149.400 17.200 ;
        RECT 149.100 16.200 149.400 16.800 ;
        RECT 144.600 15.900 145.700 16.200 ;
        RECT 148.300 15.900 148.800 16.200 ;
        RECT 149.100 15.900 149.800 16.200 ;
        RECT 142.100 15.300 144.200 15.600 ;
        RECT 142.100 15.200 142.500 15.300 ;
        RECT 143.800 15.100 144.200 15.300 ;
        RECT 145.400 15.600 145.700 15.900 ;
        RECT 145.400 15.200 146.000 15.600 ;
        RECT 144.600 15.100 145.000 15.200 ;
        RECT 142.900 14.900 143.300 15.000 ;
        RECT 141.400 14.600 143.300 14.900 ;
        RECT 143.800 14.800 145.000 15.100 ;
        RECT 141.400 14.500 141.800 14.600 ;
        RECT 133.800 14.100 134.600 14.200 ;
        RECT 132.900 13.800 134.600 14.100 ;
        RECT 135.400 13.900 140.900 14.200 ;
        RECT 135.400 13.800 136.200 13.900 ;
        RECT 132.900 13.600 133.200 13.800 ;
        RECT 132.200 13.300 133.200 13.600 ;
        RECT 133.500 13.400 133.900 13.500 ;
        RECT 132.200 13.200 133.000 13.300 ;
        RECT 133.500 13.100 134.600 13.400 ;
        RECT 131.600 11.100 132.400 12.900 ;
        RECT 134.200 11.100 134.600 13.100 ;
        RECT 135.000 11.100 135.400 13.500 ;
        RECT 137.500 12.800 137.800 13.900 ;
        RECT 140.300 13.800 140.700 13.900 ;
        RECT 143.800 13.600 144.200 14.800 ;
        RECT 144.600 14.400 145.000 14.800 ;
        RECT 145.400 13.700 145.700 15.200 ;
        RECT 147.000 15.100 147.400 15.200 ;
        RECT 147.800 15.100 148.200 15.200 ;
        RECT 147.000 14.800 148.200 15.100 ;
        RECT 147.800 14.400 148.200 14.800 ;
        RECT 148.500 14.200 148.800 15.900 ;
        RECT 149.400 15.800 149.800 15.900 ;
        RECT 147.000 14.100 147.400 14.200 ;
        RECT 147.000 13.800 147.800 14.100 ;
        RECT 148.500 13.800 149.800 14.200 ;
        RECT 142.300 13.300 144.200 13.600 ;
        RECT 142.300 13.200 142.700 13.300 ;
        RECT 136.600 12.100 137.000 12.500 ;
        RECT 137.400 12.400 137.800 12.800 ;
        RECT 138.300 12.700 138.700 12.800 ;
        RECT 138.300 12.400 139.700 12.700 ;
        RECT 139.400 12.100 139.700 12.400 ;
        RECT 141.400 12.100 141.800 12.500 ;
        RECT 136.600 11.800 137.600 12.100 ;
        RECT 137.200 11.100 137.600 11.800 ;
        RECT 139.400 11.100 139.800 12.100 ;
        RECT 141.400 11.800 142.100 12.100 ;
        RECT 141.500 11.100 142.100 11.800 ;
        RECT 143.800 11.100 144.200 13.300 ;
        RECT 144.600 13.400 145.700 13.700 ;
        RECT 147.400 13.600 147.800 13.800 ;
        RECT 144.600 11.100 145.000 13.400 ;
        RECT 147.100 13.100 148.900 13.300 ;
        RECT 149.400 13.100 149.700 13.800 ;
        RECT 147.000 13.000 149.000 13.100 ;
        RECT 147.000 11.100 147.400 13.000 ;
        RECT 148.600 11.100 149.000 13.000 ;
        RECT 149.400 11.100 149.800 13.100 ;
        RECT 0.600 7.900 1.000 9.900 ;
        RECT 2.800 9.200 3.600 9.900 ;
        RECT 2.800 8.800 4.200 9.200 ;
        RECT 2.800 8.100 3.600 8.800 ;
        RECT 0.600 7.600 1.900 7.900 ;
        RECT 1.500 7.500 1.900 7.600 ;
        RECT 2.200 7.400 3.000 7.800 ;
        RECT 3.300 7.100 3.600 8.100 ;
        RECT 5.400 7.900 5.800 9.900 ;
        RECT 7.500 8.200 7.900 9.900 ;
        RECT 3.900 7.400 4.300 7.800 ;
        RECT 4.600 7.600 5.800 7.900 ;
        RECT 7.000 7.900 7.900 8.200 ;
        RECT 8.600 7.900 9.000 9.900 ;
        RECT 9.400 8.000 9.800 9.900 ;
        RECT 11.000 8.000 11.400 9.900 ;
        RECT 9.400 7.900 11.400 8.000 ;
        RECT 11.800 7.900 12.200 9.900 ;
        RECT 14.000 9.200 14.800 9.900 ;
        RECT 14.000 8.800 15.400 9.200 ;
        RECT 14.000 8.100 14.800 8.800 ;
        RECT 4.600 7.500 5.000 7.600 ;
        RECT 3.100 6.800 3.600 7.100 ;
        RECT 4.000 7.200 4.300 7.400 ;
        RECT 4.000 6.800 4.400 7.200 ;
        RECT 6.200 6.800 6.600 7.600 ;
        RECT 3.100 6.200 3.400 6.800 ;
        RECT 1.700 6.100 2.100 6.200 ;
        RECT 1.700 5.800 2.500 6.100 ;
        RECT 3.000 5.800 3.400 6.200 ;
        RECT 2.100 5.700 2.500 5.800 ;
        RECT 3.100 5.100 3.400 5.800 ;
        RECT 6.200 5.100 6.600 5.200 ;
        RECT 7.000 5.100 7.400 7.900 ;
        RECT 8.700 7.200 9.000 7.900 ;
        RECT 9.500 7.700 11.300 7.900 ;
        RECT 11.800 7.600 13.000 7.900 ;
        RECT 12.600 7.500 13.000 7.600 ;
        RECT 13.300 7.400 13.700 7.800 ;
        RECT 10.600 7.200 11.000 7.400 ;
        RECT 13.300 7.200 13.600 7.400 ;
        RECT 8.600 6.800 9.900 7.200 ;
        RECT 10.600 6.900 11.400 7.200 ;
        RECT 11.000 6.800 11.400 6.900 ;
        RECT 11.800 6.800 12.600 7.200 ;
        RECT 13.200 6.800 13.600 7.200 ;
        RECT 14.000 7.100 14.300 8.100 ;
        RECT 16.600 7.900 17.000 9.900 ;
        RECT 17.400 7.900 17.800 9.900 ;
        RECT 18.200 8.000 18.600 9.900 ;
        RECT 19.800 8.000 20.200 9.900 ;
        RECT 18.200 7.900 20.200 8.000 ;
        RECT 14.600 7.400 15.400 7.800 ;
        RECT 15.700 7.600 17.000 7.900 ;
        RECT 15.700 7.500 16.100 7.600 ;
        RECT 17.500 7.200 17.800 7.900 ;
        RECT 18.300 7.700 20.100 7.900 ;
        RECT 19.400 7.200 19.800 7.400 ;
        RECT 16.200 7.100 17.000 7.200 ;
        RECT 17.400 7.100 18.700 7.200 ;
        RECT 14.000 6.800 14.500 7.100 ;
        RECT 15.900 7.000 18.700 7.100 ;
        RECT 0.600 4.800 1.900 5.100 ;
        RECT 0.600 1.100 1.000 4.800 ;
        RECT 1.500 4.700 1.900 4.800 ;
        RECT 2.800 1.100 3.600 5.100 ;
        RECT 4.600 4.800 5.800 5.100 ;
        RECT 6.200 4.800 7.400 5.100 ;
        RECT 4.600 4.700 5.000 4.800 ;
        RECT 5.400 1.100 5.800 4.800 ;
        RECT 7.000 1.100 7.400 4.800 ;
        RECT 7.800 4.400 8.200 5.200 ;
        RECT 8.600 5.100 9.000 5.200 ;
        RECT 9.600 5.100 9.900 6.800 ;
        RECT 14.200 6.200 14.500 6.800 ;
        RECT 14.800 6.800 18.700 7.000 ;
        RECT 19.400 7.100 20.200 7.200 ;
        RECT 20.600 7.100 21.000 9.900 ;
        RECT 22.200 7.900 22.600 9.900 ;
        RECT 24.400 9.200 25.200 9.900 ;
        RECT 24.400 8.800 25.800 9.200 ;
        RECT 24.400 8.100 25.200 8.800 ;
        RECT 22.200 7.600 23.300 7.900 ;
        RECT 22.900 7.500 23.300 7.600 ;
        RECT 19.400 6.900 21.000 7.100 ;
        RECT 19.800 6.800 21.000 6.900 ;
        RECT 14.800 6.700 16.200 6.800 ;
        RECT 14.800 6.600 15.200 6.700 ;
        RECT 14.200 5.800 14.600 6.200 ;
        RECT 15.500 6.100 15.900 6.200 ;
        RECT 15.100 5.800 15.900 6.100 ;
        RECT 14.200 5.100 14.500 5.800 ;
        RECT 15.100 5.700 15.500 5.800 ;
        RECT 17.400 5.100 17.800 5.200 ;
        RECT 18.400 5.100 18.700 6.800 ;
        RECT 8.600 4.800 9.300 5.100 ;
        RECT 9.600 4.800 10.100 5.100 ;
        RECT 9.000 4.200 9.300 4.800 ;
        RECT 9.000 3.800 9.400 4.200 ;
        RECT 9.700 1.100 10.100 4.800 ;
        RECT 11.800 4.800 13.000 5.100 ;
        RECT 11.800 1.100 12.200 4.800 ;
        RECT 12.600 4.700 13.000 4.800 ;
        RECT 14.000 1.100 14.800 5.100 ;
        RECT 15.700 4.800 17.000 5.100 ;
        RECT 17.400 4.800 18.100 5.100 ;
        RECT 18.400 4.800 18.900 5.100 ;
        RECT 15.700 4.700 16.100 4.800 ;
        RECT 16.600 1.100 17.000 4.800 ;
        RECT 17.800 4.200 18.100 4.800 ;
        RECT 17.800 3.800 18.200 4.200 ;
        RECT 18.500 1.100 18.900 4.800 ;
        RECT 20.600 1.100 21.000 6.800 ;
        RECT 24.200 6.700 24.600 7.100 ;
        RECT 24.200 6.400 24.500 6.700 ;
        RECT 23.200 6.100 24.500 6.400 ;
        RECT 24.900 6.400 25.200 8.100 ;
        RECT 27.000 7.900 27.400 9.900 ;
        RECT 27.800 7.900 28.200 9.900 ;
        RECT 28.600 8.000 29.000 9.900 ;
        RECT 30.200 8.000 30.600 9.900 ;
        RECT 28.600 7.900 30.600 8.000 ;
        RECT 31.800 8.800 32.200 9.900 ;
        RECT 26.200 7.600 27.400 7.900 ;
        RECT 26.200 7.500 26.600 7.600 ;
        RECT 27.900 7.200 28.200 7.900 ;
        RECT 28.700 7.700 30.500 7.900 ;
        RECT 31.800 7.200 32.100 8.800 ;
        RECT 27.800 6.800 29.100 7.200 ;
        RECT 24.900 6.200 25.400 6.400 ;
        RECT 24.900 6.100 25.800 6.200 ;
        RECT 23.200 6.000 23.600 6.100 ;
        RECT 25.100 5.800 28.100 6.100 ;
        RECT 24.300 5.700 24.700 5.800 ;
        RECT 23.000 5.400 24.700 5.700 ;
        RECT 23.000 5.100 23.300 5.400 ;
        RECT 25.100 5.100 25.400 5.800 ;
        RECT 27.800 5.200 28.100 5.800 ;
        RECT 27.800 5.100 28.200 5.200 ;
        RECT 28.800 5.100 29.100 6.800 ;
        RECT 31.800 6.800 32.200 7.200 ;
        RECT 32.600 6.800 33.000 7.200 ;
        RECT 29.400 6.100 29.800 6.600 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 29.400 5.800 31.400 6.100 ;
        RECT 31.000 5.400 31.400 5.800 ;
        RECT 31.800 5.100 32.100 6.800 ;
        RECT 32.600 6.100 32.900 6.800 ;
        RECT 33.400 6.100 33.800 9.900 ;
        RECT 35.000 7.900 35.400 9.900 ;
        RECT 37.200 9.200 38.000 9.900 ;
        RECT 36.600 8.800 38.000 9.200 ;
        RECT 37.200 8.100 38.000 8.800 ;
        RECT 35.000 7.600 36.300 7.900 ;
        RECT 35.900 7.500 36.300 7.600 ;
        RECT 36.600 7.400 37.400 7.800 ;
        RECT 37.700 7.100 38.000 8.100 ;
        RECT 39.800 7.900 40.200 9.900 ;
        RECT 38.300 7.400 38.700 7.800 ;
        RECT 39.000 7.600 40.200 7.900 ;
        RECT 39.000 7.500 39.400 7.600 ;
        RECT 40.600 7.500 41.000 9.900 ;
        RECT 42.800 9.200 43.200 9.900 ;
        RECT 42.200 8.900 43.200 9.200 ;
        RECT 45.000 8.900 45.400 9.900 ;
        RECT 47.100 9.200 47.700 9.900 ;
        RECT 47.000 8.900 47.700 9.200 ;
        RECT 49.400 9.100 49.800 9.900 ;
        RECT 51.000 9.100 51.400 9.200 ;
        RECT 42.200 8.500 42.600 8.900 ;
        RECT 45.000 8.600 45.300 8.900 ;
        RECT 43.000 8.200 43.400 8.600 ;
        RECT 43.900 8.300 45.300 8.600 ;
        RECT 47.000 8.500 47.400 8.900 ;
        RECT 49.400 8.800 51.400 9.100 ;
        RECT 43.900 8.200 44.300 8.300 ;
        RECT 37.500 6.800 38.000 7.100 ;
        RECT 38.400 7.200 38.700 7.400 ;
        RECT 38.400 6.800 38.800 7.200 ;
        RECT 41.000 7.100 41.800 7.200 ;
        RECT 43.100 7.100 43.400 8.200 ;
        RECT 47.900 7.700 48.300 7.800 ;
        RECT 49.400 7.700 49.800 8.800 ;
        RECT 47.900 7.400 49.800 7.700 ;
        RECT 51.800 7.500 52.200 9.900 ;
        RECT 54.000 9.200 54.400 9.900 ;
        RECT 53.400 8.900 54.400 9.200 ;
        RECT 56.200 8.900 56.600 9.900 ;
        RECT 58.300 9.200 58.900 9.900 ;
        RECT 58.200 8.900 58.900 9.200 ;
        RECT 53.400 8.500 53.800 8.900 ;
        RECT 56.200 8.600 56.500 8.900 ;
        RECT 54.200 7.800 54.600 8.600 ;
        RECT 55.100 8.300 56.500 8.600 ;
        RECT 58.200 8.500 58.600 8.900 ;
        RECT 55.100 8.200 55.500 8.300 ;
        RECT 44.600 7.100 45.000 7.200 ;
        RECT 45.900 7.100 46.300 7.200 ;
        RECT 41.000 6.800 46.500 7.100 ;
        RECT 37.500 6.200 37.800 6.800 ;
        RECT 42.500 6.700 42.900 6.800 ;
        RECT 32.600 5.800 33.800 6.100 ;
        RECT 36.100 6.100 36.500 6.200 ;
        RECT 36.100 5.800 36.900 6.100 ;
        RECT 37.400 5.800 37.800 6.200 ;
        RECT 22.200 4.800 23.300 5.100 ;
        RECT 22.200 1.100 22.600 4.800 ;
        RECT 22.900 4.700 23.300 4.800 ;
        RECT 24.400 4.800 25.400 5.100 ;
        RECT 26.200 4.800 27.400 5.100 ;
        RECT 27.800 4.800 28.500 5.100 ;
        RECT 28.800 4.800 29.300 5.100 ;
        RECT 24.400 1.100 25.200 4.800 ;
        RECT 26.200 4.700 26.600 4.800 ;
        RECT 27.000 1.100 27.400 4.800 ;
        RECT 28.200 4.200 28.500 4.800 ;
        RECT 28.200 3.800 28.600 4.200 ;
        RECT 28.900 1.100 29.300 4.800 ;
        RECT 31.300 4.700 32.200 5.100 ;
        RECT 31.300 1.100 31.700 4.700 ;
        RECT 33.400 1.100 33.800 5.800 ;
        RECT 36.500 5.700 36.900 5.800 ;
        RECT 37.500 5.100 37.800 5.800 ;
        RECT 40.600 5.500 43.400 5.600 ;
        RECT 40.600 5.400 43.500 5.500 ;
        RECT 40.600 5.300 45.500 5.400 ;
        RECT 35.000 4.800 36.300 5.100 ;
        RECT 35.000 1.100 35.400 4.800 ;
        RECT 35.900 4.700 36.300 4.800 ;
        RECT 37.200 1.100 38.000 5.100 ;
        RECT 39.000 4.800 40.200 5.100 ;
        RECT 39.000 4.700 39.400 4.800 ;
        RECT 39.800 1.100 40.200 4.800 ;
        RECT 40.600 1.100 41.000 5.300 ;
        RECT 43.100 5.100 45.500 5.300 ;
        RECT 42.200 4.500 44.900 4.800 ;
        RECT 42.200 4.400 42.600 4.500 ;
        RECT 44.500 4.400 44.900 4.500 ;
        RECT 45.200 4.500 45.500 5.100 ;
        RECT 46.200 5.200 46.500 6.800 ;
        RECT 47.000 6.400 47.400 6.500 ;
        RECT 47.000 6.100 48.900 6.400 ;
        RECT 48.500 6.000 48.900 6.100 ;
        RECT 47.700 5.700 48.100 5.800 ;
        RECT 49.400 5.700 49.800 7.400 ;
        RECT 52.200 7.100 53.000 7.200 ;
        RECT 54.300 7.100 54.600 7.800 ;
        RECT 59.100 7.700 59.500 7.800 ;
        RECT 60.600 7.700 61.000 9.900 ;
        RECT 59.100 7.400 61.000 7.700 ;
        RECT 63.000 7.600 63.400 9.900 ;
        RECT 57.100 7.100 57.500 7.200 ;
        RECT 52.200 6.800 57.700 7.100 ;
        RECT 53.700 6.700 54.100 6.800 ;
        RECT 47.700 5.400 49.800 5.700 ;
        RECT 46.200 4.900 47.400 5.200 ;
        RECT 45.900 4.500 46.300 4.600 ;
        RECT 45.200 4.200 46.300 4.500 ;
        RECT 47.100 4.400 47.400 4.900 ;
        RECT 47.100 4.000 47.800 4.400 ;
        RECT 43.900 3.700 44.300 3.800 ;
        RECT 45.300 3.700 45.700 3.800 ;
        RECT 42.200 3.100 42.600 3.500 ;
        RECT 43.900 3.400 45.700 3.700 ;
        RECT 45.000 3.100 45.300 3.400 ;
        RECT 47.000 3.100 47.400 3.500 ;
        RECT 42.200 2.800 43.200 3.100 ;
        RECT 42.800 1.100 43.200 2.800 ;
        RECT 45.000 1.100 45.400 3.100 ;
        RECT 47.100 1.100 47.700 3.100 ;
        RECT 49.400 1.100 49.800 5.400 ;
        RECT 51.800 5.500 54.600 5.600 ;
        RECT 51.800 5.400 54.700 5.500 ;
        RECT 51.800 5.300 56.700 5.400 ;
        RECT 51.800 1.100 52.200 5.300 ;
        RECT 54.300 5.100 56.700 5.300 ;
        RECT 53.400 4.500 56.100 4.800 ;
        RECT 53.400 4.400 53.800 4.500 ;
        RECT 55.700 4.400 56.100 4.500 ;
        RECT 56.400 4.500 56.700 5.100 ;
        RECT 57.400 5.200 57.700 6.800 ;
        RECT 58.200 6.400 58.600 6.500 ;
        RECT 58.200 6.100 60.100 6.400 ;
        RECT 59.700 6.000 60.100 6.100 ;
        RECT 58.900 5.700 59.300 5.800 ;
        RECT 60.600 5.700 61.000 7.400 ;
        RECT 62.300 7.300 63.400 7.600 ;
        RECT 63.800 7.700 64.200 9.900 ;
        RECT 65.900 9.200 66.500 9.900 ;
        RECT 65.900 8.900 66.600 9.200 ;
        RECT 68.200 8.900 68.600 9.900 ;
        RECT 70.400 9.200 70.800 9.900 ;
        RECT 70.400 8.900 71.400 9.200 ;
        RECT 66.200 8.500 66.600 8.900 ;
        RECT 68.300 8.600 68.600 8.900 ;
        RECT 68.300 8.300 69.700 8.600 ;
        RECT 69.300 8.200 69.700 8.300 ;
        RECT 70.200 8.200 70.600 8.600 ;
        RECT 71.000 8.500 71.400 8.900 ;
        RECT 65.300 7.700 65.700 7.800 ;
        RECT 63.800 7.400 65.700 7.700 ;
        RECT 62.300 5.800 62.600 7.300 ;
        RECT 63.000 6.100 63.400 6.600 ;
        RECT 63.800 6.100 64.200 7.400 ;
        RECT 67.300 7.100 67.700 7.200 ;
        RECT 70.200 7.100 70.500 8.200 ;
        RECT 72.600 7.500 73.000 9.900 ;
        RECT 75.000 7.600 75.400 9.900 ;
        RECT 74.300 7.300 75.400 7.600 ;
        RECT 75.800 7.700 76.200 9.900 ;
        RECT 77.900 9.200 78.500 9.900 ;
        RECT 77.900 8.900 78.600 9.200 ;
        RECT 80.200 8.900 80.600 9.900 ;
        RECT 82.400 9.200 82.800 9.900 ;
        RECT 82.400 8.900 83.400 9.200 ;
        RECT 78.200 8.500 78.600 8.900 ;
        RECT 80.300 8.600 80.600 8.900 ;
        RECT 80.300 8.300 81.700 8.600 ;
        RECT 81.300 8.200 81.700 8.300 ;
        RECT 82.200 8.200 82.600 8.600 ;
        RECT 83.000 8.500 83.400 8.900 ;
        RECT 77.300 7.700 77.700 7.800 ;
        RECT 75.800 7.400 77.700 7.700 ;
        RECT 71.800 7.100 72.600 7.200 ;
        RECT 67.100 6.800 72.600 7.100 ;
        RECT 66.200 6.400 66.600 6.500 ;
        RECT 63.000 5.800 64.200 6.100 ;
        RECT 64.700 6.100 66.600 6.400 ;
        RECT 64.700 6.000 65.100 6.100 ;
        RECT 58.900 5.400 61.000 5.700 ;
        RECT 62.000 5.400 62.600 5.800 ;
        RECT 57.400 4.900 58.600 5.200 ;
        RECT 57.100 4.500 57.500 4.600 ;
        RECT 56.400 4.200 57.500 4.500 ;
        RECT 58.300 4.400 58.600 4.900 ;
        RECT 58.300 4.000 59.000 4.400 ;
        RECT 55.100 3.700 55.500 3.800 ;
        RECT 56.500 3.700 56.900 3.800 ;
        RECT 53.400 3.100 53.800 3.500 ;
        RECT 55.100 3.400 56.900 3.700 ;
        RECT 56.200 3.100 56.500 3.400 ;
        RECT 58.200 3.100 58.600 3.500 ;
        RECT 53.400 2.800 54.400 3.100 ;
        RECT 54.000 1.100 54.400 2.800 ;
        RECT 56.200 1.100 56.600 3.100 ;
        RECT 58.300 1.100 58.900 3.100 ;
        RECT 60.600 1.100 61.000 5.400 ;
        RECT 62.300 5.100 62.600 5.400 ;
        RECT 63.800 5.700 64.200 5.800 ;
        RECT 65.500 5.700 65.900 5.800 ;
        RECT 63.800 5.400 65.900 5.700 ;
        RECT 62.300 4.800 63.400 5.100 ;
        RECT 63.000 1.100 63.400 4.800 ;
        RECT 63.800 1.100 64.200 5.400 ;
        RECT 67.100 5.200 67.400 6.800 ;
        RECT 70.700 6.700 71.100 6.800 ;
        RECT 70.200 6.200 70.600 6.300 ;
        RECT 71.500 6.200 71.900 6.300 ;
        RECT 69.400 5.900 71.900 6.200 ;
        RECT 69.400 5.800 69.800 5.900 ;
        RECT 74.300 5.800 74.600 7.300 ;
        RECT 75.000 6.100 75.400 6.600 ;
        RECT 75.800 6.100 76.200 7.400 ;
        RECT 79.300 7.100 79.700 7.200 ;
        RECT 80.600 7.100 81.000 7.200 ;
        RECT 82.200 7.100 82.500 8.200 ;
        RECT 84.600 7.500 85.000 9.900 ;
        RECT 85.400 7.500 85.800 9.900 ;
        RECT 87.600 9.200 88.000 9.900 ;
        RECT 87.000 8.900 88.000 9.200 ;
        RECT 89.800 8.900 90.200 9.900 ;
        RECT 91.900 9.200 92.500 9.900 ;
        RECT 91.800 8.900 92.500 9.200 ;
        RECT 87.000 8.500 87.400 8.900 ;
        RECT 89.800 8.600 90.100 8.900 ;
        RECT 87.800 8.200 88.200 8.600 ;
        RECT 88.700 8.300 90.100 8.600 ;
        RECT 91.800 8.500 92.200 8.900 ;
        RECT 88.700 8.200 89.100 8.300 ;
        RECT 83.800 7.100 84.600 7.200 ;
        RECT 85.800 7.100 86.600 7.200 ;
        RECT 87.900 7.100 88.200 8.200 ;
        RECT 91.000 7.800 91.400 8.200 ;
        RECT 91.000 7.200 91.300 7.800 ;
        RECT 92.700 7.700 93.100 7.800 ;
        RECT 94.200 7.700 94.600 9.900 ;
        RECT 92.700 7.400 94.600 7.700 ;
        RECT 90.700 7.100 91.300 7.200 ;
        RECT 79.100 6.800 91.300 7.100 ;
        RECT 78.200 6.400 78.600 6.500 ;
        RECT 75.000 5.800 76.200 6.100 ;
        RECT 76.700 6.100 78.600 6.400 ;
        RECT 76.700 6.000 77.100 6.100 ;
        RECT 70.200 5.500 73.000 5.600 ;
        RECT 70.100 5.400 73.000 5.500 ;
        RECT 74.000 5.400 74.600 5.800 ;
        RECT 66.200 4.900 67.400 5.200 ;
        RECT 68.100 5.300 73.000 5.400 ;
        RECT 68.100 5.100 70.500 5.300 ;
        RECT 66.200 4.400 66.500 4.900 ;
        RECT 65.800 4.000 66.500 4.400 ;
        RECT 67.300 4.500 67.700 4.600 ;
        RECT 68.100 4.500 68.400 5.100 ;
        RECT 67.300 4.200 68.400 4.500 ;
        RECT 68.700 4.500 71.400 4.800 ;
        RECT 68.700 4.400 69.100 4.500 ;
        RECT 71.000 4.400 71.400 4.500 ;
        RECT 67.900 3.700 68.300 3.800 ;
        RECT 69.300 3.700 69.700 3.800 ;
        RECT 66.200 3.100 66.600 3.500 ;
        RECT 67.900 3.400 69.700 3.700 ;
        RECT 68.300 3.100 68.600 3.400 ;
        RECT 71.000 3.100 71.400 3.500 ;
        RECT 65.900 1.100 66.500 3.100 ;
        RECT 68.200 1.100 68.600 3.100 ;
        RECT 70.400 2.800 71.400 3.100 ;
        RECT 70.400 1.100 70.800 2.800 ;
        RECT 72.600 1.100 73.000 5.300 ;
        RECT 74.300 5.100 74.600 5.400 ;
        RECT 75.800 5.700 76.200 5.800 ;
        RECT 77.500 5.700 77.900 5.800 ;
        RECT 75.800 5.400 77.900 5.700 ;
        RECT 74.300 4.800 75.400 5.100 ;
        RECT 75.000 1.100 75.400 4.800 ;
        RECT 75.800 1.100 76.200 5.400 ;
        RECT 79.100 5.200 79.400 6.800 ;
        RECT 82.700 6.700 83.100 6.800 ;
        RECT 87.300 6.700 87.700 6.800 ;
        RECT 82.200 6.200 82.600 6.300 ;
        RECT 83.500 6.200 83.900 6.300 ;
        RECT 81.400 5.900 83.900 6.200 ;
        RECT 86.500 6.200 86.900 6.300 ;
        RECT 87.800 6.200 88.200 6.300 ;
        RECT 86.500 5.900 89.000 6.200 ;
        RECT 81.400 5.800 81.800 5.900 ;
        RECT 88.600 5.800 89.000 5.900 ;
        RECT 82.200 5.500 85.000 5.600 ;
        RECT 82.100 5.400 85.000 5.500 ;
        RECT 78.200 4.900 79.400 5.200 ;
        RECT 80.100 5.300 85.000 5.400 ;
        RECT 80.100 5.100 82.500 5.300 ;
        RECT 78.200 4.400 78.500 4.900 ;
        RECT 77.800 4.000 78.500 4.400 ;
        RECT 79.300 4.500 79.700 4.600 ;
        RECT 80.100 4.500 80.400 5.100 ;
        RECT 79.300 4.200 80.400 4.500 ;
        RECT 80.700 4.500 83.400 4.800 ;
        RECT 80.700 4.400 81.100 4.500 ;
        RECT 83.000 4.400 83.400 4.500 ;
        RECT 79.900 3.700 80.300 3.800 ;
        RECT 81.300 3.700 81.700 3.800 ;
        RECT 78.200 3.100 78.600 3.500 ;
        RECT 79.900 3.400 81.700 3.700 ;
        RECT 80.300 3.100 80.600 3.400 ;
        RECT 83.000 3.100 83.400 3.500 ;
        RECT 77.900 1.100 78.500 3.100 ;
        RECT 80.200 1.100 80.600 3.100 ;
        RECT 82.400 2.800 83.400 3.100 ;
        RECT 82.400 1.100 82.800 2.800 ;
        RECT 84.600 1.100 85.000 5.300 ;
        RECT 85.400 5.500 88.200 5.600 ;
        RECT 85.400 5.400 88.300 5.500 ;
        RECT 85.400 5.300 90.300 5.400 ;
        RECT 85.400 1.100 85.800 5.300 ;
        RECT 87.900 5.100 90.300 5.300 ;
        RECT 87.000 4.500 89.700 4.800 ;
        RECT 87.000 4.400 87.400 4.500 ;
        RECT 89.300 4.400 89.700 4.500 ;
        RECT 90.000 4.500 90.300 5.100 ;
        RECT 91.000 5.200 91.300 6.800 ;
        RECT 91.800 6.400 92.200 6.500 ;
        RECT 91.800 6.100 93.700 6.400 ;
        RECT 93.300 6.000 93.700 6.100 ;
        RECT 94.200 6.100 94.600 7.400 ;
        RECT 95.000 7.600 95.400 9.900 ;
        RECT 95.000 7.300 96.100 7.600 ;
        RECT 99.000 7.500 99.400 9.900 ;
        RECT 101.200 9.200 101.600 9.900 ;
        RECT 100.600 8.900 101.600 9.200 ;
        RECT 103.400 8.900 103.800 9.900 ;
        RECT 105.500 9.200 106.100 9.900 ;
        RECT 105.400 8.900 106.100 9.200 ;
        RECT 100.600 8.500 101.000 8.900 ;
        RECT 103.400 8.600 103.700 8.900 ;
        RECT 101.400 8.200 101.800 8.600 ;
        RECT 102.300 8.300 103.700 8.600 ;
        RECT 105.400 8.500 105.800 8.900 ;
        RECT 102.300 8.200 102.700 8.300 ;
        RECT 95.000 6.100 95.400 6.600 ;
        RECT 94.200 5.800 95.400 6.100 ;
        RECT 95.800 5.800 96.100 7.300 ;
        RECT 99.400 7.100 100.200 7.200 ;
        RECT 101.500 7.100 101.800 8.200 ;
        RECT 106.300 7.700 106.700 7.800 ;
        RECT 107.800 7.700 108.200 9.900 ;
        RECT 106.300 7.400 108.200 7.700 ;
        RECT 104.300 7.100 104.700 7.200 ;
        RECT 99.400 6.800 104.900 7.100 ;
        RECT 100.900 6.700 101.300 6.800 ;
        RECT 100.100 6.200 100.500 6.300 ;
        RECT 101.400 6.200 101.800 6.300 ;
        RECT 100.100 5.900 102.600 6.200 ;
        RECT 102.200 5.800 102.600 5.900 ;
        RECT 92.500 5.700 92.900 5.800 ;
        RECT 94.200 5.700 94.600 5.800 ;
        RECT 92.500 5.400 94.600 5.700 ;
        RECT 91.000 4.900 92.200 5.200 ;
        RECT 90.700 4.500 91.100 4.600 ;
        RECT 90.000 4.200 91.100 4.500 ;
        RECT 91.900 4.400 92.200 4.900 ;
        RECT 91.900 4.000 92.600 4.400 ;
        RECT 88.700 3.700 89.100 3.800 ;
        RECT 90.100 3.700 90.500 3.800 ;
        RECT 87.000 3.100 87.400 3.500 ;
        RECT 88.700 3.400 90.500 3.700 ;
        RECT 89.800 3.100 90.100 3.400 ;
        RECT 91.800 3.100 92.200 3.500 ;
        RECT 87.000 2.800 88.000 3.100 ;
        RECT 87.600 1.100 88.000 2.800 ;
        RECT 89.800 1.100 90.200 3.100 ;
        RECT 91.900 1.100 92.500 3.100 ;
        RECT 94.200 1.100 94.600 5.400 ;
        RECT 95.800 5.400 96.400 5.800 ;
        RECT 99.000 5.500 101.800 5.600 ;
        RECT 99.000 5.400 101.900 5.500 ;
        RECT 95.800 5.100 96.100 5.400 ;
        RECT 95.000 4.800 96.100 5.100 ;
        RECT 99.000 5.300 103.900 5.400 ;
        RECT 95.000 1.100 95.400 4.800 ;
        RECT 99.000 1.100 99.400 5.300 ;
        RECT 101.500 5.100 103.900 5.300 ;
        RECT 100.600 4.500 103.300 4.800 ;
        RECT 100.600 4.400 101.000 4.500 ;
        RECT 102.900 4.400 103.300 4.500 ;
        RECT 103.600 4.500 103.900 5.100 ;
        RECT 104.600 5.200 104.900 6.800 ;
        RECT 105.400 6.400 105.800 6.500 ;
        RECT 105.400 6.100 107.300 6.400 ;
        RECT 106.900 6.000 107.300 6.100 ;
        RECT 107.800 6.100 108.200 7.400 ;
        RECT 108.600 7.600 109.000 9.900 ;
        RECT 108.600 7.300 109.700 7.600 ;
        RECT 111.000 7.500 111.400 9.900 ;
        RECT 113.200 9.200 113.600 9.900 ;
        RECT 112.600 8.900 113.600 9.200 ;
        RECT 115.400 8.900 115.800 9.900 ;
        RECT 117.500 9.200 118.100 9.900 ;
        RECT 117.400 8.900 118.100 9.200 ;
        RECT 112.600 8.500 113.000 8.900 ;
        RECT 115.400 8.600 115.700 8.900 ;
        RECT 113.400 8.200 113.800 8.600 ;
        RECT 114.300 8.300 115.700 8.600 ;
        RECT 117.400 8.500 117.800 8.900 ;
        RECT 114.300 8.200 114.700 8.300 ;
        RECT 108.600 6.100 109.000 6.600 ;
        RECT 107.800 5.800 109.000 6.100 ;
        RECT 109.400 5.800 109.700 7.300 ;
        RECT 111.400 7.100 112.200 7.200 ;
        RECT 113.500 7.100 113.800 8.200 ;
        RECT 118.300 7.700 118.700 7.800 ;
        RECT 119.800 7.700 120.200 9.900 ;
        RECT 118.300 7.400 120.200 7.700 ;
        RECT 116.300 7.100 116.700 7.200 ;
        RECT 111.400 6.800 116.900 7.100 ;
        RECT 112.900 6.700 113.300 6.800 ;
        RECT 112.100 6.200 112.500 6.300 ;
        RECT 113.400 6.200 113.800 6.300 ;
        RECT 112.100 5.900 114.600 6.200 ;
        RECT 114.200 5.800 114.600 5.900 ;
        RECT 106.100 5.700 106.500 5.800 ;
        RECT 107.800 5.700 108.200 5.800 ;
        RECT 106.100 5.400 108.200 5.700 ;
        RECT 104.600 4.900 105.800 5.200 ;
        RECT 104.300 4.500 104.700 4.600 ;
        RECT 103.600 4.200 104.700 4.500 ;
        RECT 105.500 4.400 105.800 4.900 ;
        RECT 105.500 4.000 106.200 4.400 ;
        RECT 102.300 3.700 102.700 3.800 ;
        RECT 103.700 3.700 104.100 3.800 ;
        RECT 100.600 3.100 101.000 3.500 ;
        RECT 102.300 3.400 104.100 3.700 ;
        RECT 103.400 3.100 103.700 3.400 ;
        RECT 105.400 3.100 105.800 3.500 ;
        RECT 100.600 2.800 101.600 3.100 ;
        RECT 101.200 1.100 101.600 2.800 ;
        RECT 103.400 1.100 103.800 3.100 ;
        RECT 105.500 1.100 106.100 3.100 ;
        RECT 107.800 1.100 108.200 5.400 ;
        RECT 109.400 5.400 110.000 5.800 ;
        RECT 111.000 5.500 113.800 5.600 ;
        RECT 111.000 5.400 113.900 5.500 ;
        RECT 109.400 5.100 109.700 5.400 ;
        RECT 108.600 4.800 109.700 5.100 ;
        RECT 111.000 5.300 115.900 5.400 ;
        RECT 108.600 1.100 109.000 4.800 ;
        RECT 111.000 1.100 111.400 5.300 ;
        RECT 113.500 5.100 115.900 5.300 ;
        RECT 112.600 4.500 115.300 4.800 ;
        RECT 112.600 4.400 113.000 4.500 ;
        RECT 114.900 4.400 115.300 4.500 ;
        RECT 115.600 4.500 115.900 5.100 ;
        RECT 116.600 5.200 116.900 6.800 ;
        RECT 117.400 6.400 117.800 6.500 ;
        RECT 117.400 6.100 119.300 6.400 ;
        RECT 118.900 6.000 119.300 6.100 ;
        RECT 119.800 6.100 120.200 7.400 ;
        RECT 120.600 7.600 121.000 9.900 ;
        RECT 120.600 7.300 121.700 7.600 ;
        RECT 123.000 7.500 123.400 9.900 ;
        RECT 125.200 9.200 125.600 9.900 ;
        RECT 124.600 8.900 125.600 9.200 ;
        RECT 127.400 8.900 127.800 9.900 ;
        RECT 129.500 9.200 130.100 9.900 ;
        RECT 129.400 8.900 130.100 9.200 ;
        RECT 124.600 8.500 125.000 8.900 ;
        RECT 127.400 8.600 127.700 8.900 ;
        RECT 125.400 8.200 125.800 8.600 ;
        RECT 126.300 8.300 127.700 8.600 ;
        RECT 129.400 8.500 129.800 8.900 ;
        RECT 126.300 8.200 126.700 8.300 ;
        RECT 120.600 6.100 121.000 6.600 ;
        RECT 119.800 5.800 121.000 6.100 ;
        RECT 121.400 5.800 121.700 7.300 ;
        RECT 123.400 7.100 124.200 7.200 ;
        RECT 125.500 7.100 125.800 8.200 ;
        RECT 130.300 7.700 130.700 7.800 ;
        RECT 131.800 7.700 132.200 9.900 ;
        RECT 130.300 7.400 132.200 7.700 ;
        RECT 128.300 7.100 128.700 7.200 ;
        RECT 123.400 6.800 128.900 7.100 ;
        RECT 124.900 6.700 125.300 6.800 ;
        RECT 124.100 6.200 124.500 6.300 ;
        RECT 125.400 6.200 125.800 6.300 ;
        RECT 124.100 5.900 126.600 6.200 ;
        RECT 126.200 5.800 126.600 5.900 ;
        RECT 118.100 5.700 118.500 5.800 ;
        RECT 119.800 5.700 120.200 5.800 ;
        RECT 118.100 5.400 120.200 5.700 ;
        RECT 116.600 4.900 117.800 5.200 ;
        RECT 116.300 4.500 116.700 4.600 ;
        RECT 115.600 4.200 116.700 4.500 ;
        RECT 117.500 4.400 117.800 4.900 ;
        RECT 117.500 4.000 118.200 4.400 ;
        RECT 114.300 3.700 114.700 3.800 ;
        RECT 115.700 3.700 116.100 3.800 ;
        RECT 112.600 3.100 113.000 3.500 ;
        RECT 114.300 3.400 116.100 3.700 ;
        RECT 115.400 3.100 115.700 3.400 ;
        RECT 117.400 3.100 117.800 3.500 ;
        RECT 112.600 2.800 113.600 3.100 ;
        RECT 113.200 1.100 113.600 2.800 ;
        RECT 115.400 1.100 115.800 3.100 ;
        RECT 117.500 1.100 118.100 3.100 ;
        RECT 119.800 1.100 120.200 5.400 ;
        RECT 121.400 5.400 122.000 5.800 ;
        RECT 123.000 5.500 125.800 5.600 ;
        RECT 123.000 5.400 125.900 5.500 ;
        RECT 121.400 5.100 121.700 5.400 ;
        RECT 120.600 4.800 121.700 5.100 ;
        RECT 123.000 5.300 127.900 5.400 ;
        RECT 120.600 1.100 121.000 4.800 ;
        RECT 123.000 1.100 123.400 5.300 ;
        RECT 125.500 5.100 127.900 5.300 ;
        RECT 124.600 4.500 127.300 4.800 ;
        RECT 124.600 4.400 125.000 4.500 ;
        RECT 126.900 4.400 127.300 4.500 ;
        RECT 127.600 4.500 127.900 5.100 ;
        RECT 128.600 5.200 128.900 6.800 ;
        RECT 129.400 6.400 129.800 6.500 ;
        RECT 129.400 6.100 131.300 6.400 ;
        RECT 130.900 6.000 131.300 6.100 ;
        RECT 131.800 6.100 132.200 7.400 ;
        RECT 132.600 7.600 133.000 9.900 ;
        RECT 132.600 7.300 133.700 7.600 ;
        RECT 135.000 7.500 135.400 9.900 ;
        RECT 137.200 9.200 137.600 9.900 ;
        RECT 136.600 8.900 137.600 9.200 ;
        RECT 139.400 8.900 139.800 9.900 ;
        RECT 141.500 9.200 142.100 9.900 ;
        RECT 141.400 8.900 142.100 9.200 ;
        RECT 136.600 8.500 137.000 8.900 ;
        RECT 139.400 8.600 139.700 8.900 ;
        RECT 137.400 8.200 137.800 8.600 ;
        RECT 138.300 8.300 139.700 8.600 ;
        RECT 141.400 8.500 141.800 8.900 ;
        RECT 138.300 8.200 138.700 8.300 ;
        RECT 132.600 6.100 133.000 6.600 ;
        RECT 131.800 5.800 133.000 6.100 ;
        RECT 133.400 5.800 133.700 7.300 ;
        RECT 135.400 7.100 136.200 7.200 ;
        RECT 137.500 7.100 137.800 8.200 ;
        RECT 142.300 7.700 142.700 7.800 ;
        RECT 143.800 7.700 144.200 9.900 ;
        RECT 142.300 7.400 144.200 7.700 ;
        RECT 140.300 7.100 140.700 7.200 ;
        RECT 135.400 6.800 140.900 7.100 ;
        RECT 136.900 6.700 137.300 6.800 ;
        RECT 136.100 6.200 136.500 6.300 ;
        RECT 136.100 5.900 138.600 6.200 ;
        RECT 138.200 5.800 138.600 5.900 ;
        RECT 130.100 5.700 130.500 5.800 ;
        RECT 131.800 5.700 132.200 5.800 ;
        RECT 130.100 5.400 132.200 5.700 ;
        RECT 128.600 4.900 129.800 5.200 ;
        RECT 128.300 4.500 128.700 4.600 ;
        RECT 127.600 4.200 128.700 4.500 ;
        RECT 129.500 4.400 129.800 4.900 ;
        RECT 129.500 4.000 130.200 4.400 ;
        RECT 126.300 3.700 126.700 3.800 ;
        RECT 127.700 3.700 128.100 3.800 ;
        RECT 124.600 3.100 125.000 3.500 ;
        RECT 126.300 3.400 128.100 3.700 ;
        RECT 127.400 3.100 127.700 3.400 ;
        RECT 129.400 3.100 129.800 3.500 ;
        RECT 124.600 2.800 125.600 3.100 ;
        RECT 125.200 1.100 125.600 2.800 ;
        RECT 127.400 1.100 127.800 3.100 ;
        RECT 129.500 1.100 130.100 3.100 ;
        RECT 131.800 1.100 132.200 5.400 ;
        RECT 133.400 5.400 134.000 5.800 ;
        RECT 135.000 5.500 137.800 5.600 ;
        RECT 135.000 5.400 137.900 5.500 ;
        RECT 133.400 5.100 133.700 5.400 ;
        RECT 132.600 4.800 133.700 5.100 ;
        RECT 135.000 5.300 139.900 5.400 ;
        RECT 132.600 1.100 133.000 4.800 ;
        RECT 135.000 1.100 135.400 5.300 ;
        RECT 137.500 5.100 139.900 5.300 ;
        RECT 136.600 4.500 139.300 4.800 ;
        RECT 136.600 4.400 137.000 4.500 ;
        RECT 138.900 4.400 139.300 4.500 ;
        RECT 139.600 4.500 139.900 5.100 ;
        RECT 140.600 5.200 140.900 6.800 ;
        RECT 141.400 6.400 141.800 6.500 ;
        RECT 141.400 6.100 143.300 6.400 ;
        RECT 142.900 6.000 143.300 6.100 ;
        RECT 143.800 6.100 144.200 7.400 ;
        RECT 144.600 7.600 145.000 9.900 ;
        RECT 147.300 9.200 147.700 9.900 ;
        RECT 147.000 8.800 147.700 9.200 ;
        RECT 147.300 8.200 147.700 8.800 ;
        RECT 147.300 7.900 148.200 8.200 ;
        RECT 144.600 7.300 145.700 7.600 ;
        RECT 144.600 6.100 145.000 6.600 ;
        RECT 143.800 5.800 145.000 6.100 ;
        RECT 145.400 5.800 145.700 7.300 ;
        RECT 142.100 5.700 142.500 5.800 ;
        RECT 143.800 5.700 144.200 5.800 ;
        RECT 142.100 5.400 144.200 5.700 ;
        RECT 140.600 4.900 141.800 5.200 ;
        RECT 140.300 4.500 140.700 4.600 ;
        RECT 139.600 4.200 140.700 4.500 ;
        RECT 141.500 4.400 141.800 4.900 ;
        RECT 141.500 4.000 142.200 4.400 ;
        RECT 138.300 3.700 138.700 3.800 ;
        RECT 139.700 3.700 140.100 3.800 ;
        RECT 136.600 3.100 137.000 3.500 ;
        RECT 138.300 3.400 140.100 3.700 ;
        RECT 139.400 3.100 139.700 3.400 ;
        RECT 141.400 3.100 141.800 3.500 ;
        RECT 136.600 2.800 137.600 3.100 ;
        RECT 137.200 1.100 137.600 2.800 ;
        RECT 139.400 1.100 139.800 3.100 ;
        RECT 141.500 1.100 142.100 3.100 ;
        RECT 143.800 1.100 144.200 5.400 ;
        RECT 145.400 5.400 146.000 5.800 ;
        RECT 145.400 5.100 145.700 5.400 ;
        RECT 144.600 4.800 145.700 5.100 ;
        RECT 144.600 1.100 145.000 4.800 ;
        RECT 147.000 4.400 147.400 5.200 ;
        RECT 147.800 1.100 148.200 7.900 ;
        RECT 148.600 6.800 149.000 7.600 ;
      LAYER via1 ;
        RECT 8.600 126.800 9.000 127.200 ;
        RECT 10.200 126.800 10.600 127.200 ;
        RECT 15.000 127.400 15.400 127.800 ;
        RECT 7.800 125.800 8.200 126.200 ;
        RECT 9.400 125.800 9.800 126.200 ;
        RECT 11.000 125.800 11.400 126.200 ;
        RECT 27.000 127.400 27.400 127.800 ;
        RECT 27.000 124.800 27.400 125.200 ;
        RECT 29.400 124.800 29.800 125.200 ;
        RECT 35.000 126.800 35.400 127.200 ;
        RECT 34.200 125.900 34.600 126.300 ;
        RECT 31.800 125.100 32.200 125.500 ;
        RECT 41.400 125.800 41.800 126.200 ;
        RECT 40.600 121.800 41.000 122.200 ;
        RECT 43.800 124.800 44.200 125.200 ;
        RECT 42.200 121.800 42.600 122.200 ;
        RECT 47.800 124.800 48.200 125.200 ;
        RECT 52.600 124.800 53.000 125.200 ;
        RECT 51.800 121.800 52.200 122.200 ;
        RECT 58.200 127.400 58.600 127.800 ;
        RECT 59.800 126.800 60.200 127.200 ;
        RECT 61.400 126.800 61.800 127.200 ;
        RECT 63.000 125.900 63.400 126.300 ;
        RECT 60.600 125.100 61.000 125.500 ;
        RECT 58.200 123.800 58.600 124.200 ;
        RECT 73.400 127.400 73.800 127.800 ;
        RECT 77.400 127.400 77.800 127.800 ;
        RECT 75.800 126.800 76.200 127.200 ;
        RECT 86.200 127.400 86.600 127.800 ;
        RECT 87.800 126.800 88.200 127.200 ;
        RECT 107.000 128.800 107.400 129.200 ;
        RECT 69.400 121.800 69.800 122.200 ;
        RECT 73.400 122.800 73.800 123.200 ;
        RECT 79.000 124.800 79.400 125.200 ;
        RECT 96.600 125.800 97.000 126.200 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 86.200 123.800 86.600 124.200 ;
        RECT 107.800 126.800 108.200 127.200 ;
        RECT 107.000 125.800 107.400 126.200 ;
        RECT 115.800 127.400 116.200 127.800 ;
        RECT 117.400 126.800 117.800 127.200 ;
        RECT 119.000 126.800 119.400 127.200 ;
        RECT 111.000 125.800 111.400 126.200 ;
        RECT 121.400 126.800 121.800 127.200 ;
        RECT 91.000 121.800 91.400 122.200 ;
        RECT 96.600 121.800 97.000 122.200 ;
        RECT 111.800 124.800 112.200 125.200 ;
        RECT 129.400 127.400 129.800 127.800 ;
        RECT 131.000 126.800 131.400 127.200 ;
        RECT 125.400 121.800 125.800 122.200 ;
        RECT 136.600 126.800 137.000 127.200 ;
        RECT 144.600 127.400 145.000 127.800 ;
        RECT 137.400 125.800 137.800 126.200 ;
        RECT 146.200 126.800 146.600 127.200 ;
        RECT 139.800 125.800 140.200 126.200 ;
        RECT 150.200 125.800 150.600 126.200 ;
        RECT 134.200 122.800 134.600 123.200 ;
        RECT 148.600 121.800 149.000 122.200 ;
        RECT 3.800 115.900 4.200 116.300 ;
        RECT 11.800 115.900 12.200 116.300 ;
        RECT 3.800 113.100 4.200 113.500 ;
        RECT 2.200 111.800 2.600 112.200 ;
        RECT 6.200 113.200 6.600 113.600 ;
        RECT 6.200 111.800 6.600 112.200 ;
        RECT 8.600 112.800 9.000 113.200 ;
        RECT 11.800 113.100 12.200 113.500 ;
        RECT 15.800 113.800 16.200 114.200 ;
        RECT 14.200 113.200 14.600 113.600 ;
        RECT 13.400 111.800 13.800 112.200 ;
        RECT 16.600 112.800 17.000 113.200 ;
        RECT 19.000 114.800 19.400 115.200 ;
        RECT 21.400 113.800 21.800 114.200 ;
        RECT 24.600 115.900 25.000 116.300 ;
        RECT 27.000 115.800 27.400 116.200 ;
        RECT 24.600 113.100 25.000 113.500 ;
        RECT 28.600 113.800 29.000 114.200 ;
        RECT 27.000 113.200 27.400 113.600 ;
        RECT 29.400 113.100 29.800 113.500 ;
        RECT 38.200 111.800 38.600 112.200 ;
        RECT 43.000 112.800 43.400 113.200 ;
        RECT 54.200 114.800 54.600 115.200 ;
        RECT 44.600 112.800 45.000 113.200 ;
        RECT 47.000 112.800 47.400 113.200 ;
        RECT 54.200 113.800 54.600 114.200 ;
        RECT 56.600 112.800 57.000 113.200 ;
        RECT 75.800 118.800 76.200 119.200 ;
        RECT 73.300 115.900 73.700 116.300 ;
        RECT 79.000 118.800 79.400 119.200 ;
        RECT 62.200 112.800 62.600 113.200 ;
        RECT 63.000 113.100 63.400 113.500 ;
        RECT 71.800 111.800 72.200 112.200 ;
        RECT 73.300 113.100 73.700 113.500 ;
        RECT 79.000 113.800 79.400 114.200 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 84.600 113.800 85.000 114.200 ;
        RECT 90.200 118.800 90.600 119.200 ;
        RECT 93.400 117.800 93.800 118.200 ;
        RECT 89.400 115.800 89.800 116.200 ;
        RECT 88.600 112.800 89.000 113.200 ;
        RECT 87.800 111.800 88.200 112.200 ;
        RECT 92.600 112.800 93.000 113.200 ;
        RECT 95.800 118.800 96.200 119.200 ;
        RECT 95.000 116.800 95.400 117.200 ;
        RECT 96.600 115.800 97.000 116.200 ;
        RECT 104.600 118.800 105.000 119.200 ;
        RECT 95.800 114.800 96.200 115.200 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 112.600 114.800 113.000 115.200 ;
        RECT 115.700 115.900 116.100 116.300 ;
        RECT 123.000 118.800 123.400 119.200 ;
        RECT 122.200 116.800 122.600 117.200 ;
        RECT 124.600 116.800 125.000 117.200 ;
        RECT 120.600 115.800 121.000 116.200 ;
        RECT 115.700 113.100 116.100 113.500 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 126.200 115.800 126.600 116.200 ;
        RECT 131.000 115.900 131.400 116.300 ;
        RECT 136.600 116.800 137.000 117.200 ;
        RECT 125.400 114.800 125.800 115.200 ;
        RECT 124.600 113.800 125.000 114.200 ;
        RECT 138.200 115.800 138.600 116.200 ;
        RECT 143.000 116.800 143.400 117.200 ;
        RECT 137.400 114.800 137.800 115.200 ;
        RECT 131.000 113.100 131.400 113.500 ;
        RECT 128.600 111.800 129.000 112.200 ;
        RECT 135.000 113.800 135.400 114.200 ;
        RECT 133.400 113.200 133.800 113.600 ;
        RECT 133.400 111.800 133.800 112.200 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 140.600 111.800 141.000 112.200 ;
        RECT 146.200 112.800 146.600 113.200 ;
        RECT 147.800 111.800 148.200 112.200 ;
        RECT 3.800 107.800 4.200 108.200 ;
        RECT 19.800 108.800 20.200 109.200 ;
        RECT 29.400 108.800 29.800 109.200 ;
        RECT 13.400 105.900 13.800 106.300 ;
        RECT 10.200 104.800 10.600 105.200 ;
        RECT 11.000 105.100 11.400 105.500 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 23.000 106.800 23.400 107.200 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 20.600 105.100 21.000 105.500 ;
        RECT 41.400 108.800 41.800 109.200 ;
        RECT 35.000 106.800 35.400 107.200 ;
        RECT 27.800 103.800 28.200 104.200 ;
        RECT 41.400 107.400 41.800 107.800 ;
        RECT 32.600 101.800 33.000 102.200 ;
        RECT 37.400 104.800 37.800 105.200 ;
        RECT 46.200 106.800 46.600 107.200 ;
        RECT 45.400 105.800 45.800 106.200 ;
        RECT 53.400 107.400 53.800 107.800 ;
        RECT 55.000 106.800 55.400 107.200 ;
        RECT 58.200 105.900 58.600 106.300 ;
        RECT 55.800 105.100 56.200 105.500 ;
        RECT 53.400 103.800 53.800 104.200 ;
        RECT 66.200 106.800 66.600 107.200 ;
        RECT 78.200 108.800 78.600 109.200 ;
        RECT 64.600 101.800 65.000 102.200 ;
        RECT 65.400 105.100 65.800 105.500 ;
        RECT 84.600 108.800 85.000 109.200 ;
        RECT 79.800 106.800 80.200 107.200 ;
        RECT 74.200 101.800 74.600 102.200 ;
        RECT 83.800 106.800 84.200 107.200 ;
        RECT 90.200 108.800 90.600 109.200 ;
        RECT 93.400 108.800 93.800 109.200 ;
        RECT 82.200 104.800 82.600 105.200 ;
        RECT 87.800 105.800 88.200 106.200 ;
        RECT 91.000 105.800 91.400 106.200 ;
        RECT 94.200 106.800 94.600 107.200 ;
        RECT 96.600 106.800 97.000 107.200 ;
        RECT 99.000 105.800 99.400 106.200 ;
        RECT 88.600 103.800 89.000 104.200 ;
        RECT 87.800 102.800 88.200 103.200 ;
        RECT 107.000 106.800 107.400 107.200 ;
        RECT 104.600 105.800 105.000 106.200 ;
        RECT 102.200 104.800 102.600 105.200 ;
        RECT 107.800 105.800 108.200 106.200 ;
        RECT 109.400 105.800 109.800 106.200 ;
        RECT 99.800 101.800 100.200 102.200 ;
        RECT 104.600 102.800 105.000 103.200 ;
        RECT 121.400 106.800 121.800 107.200 ;
        RECT 115.000 105.800 115.400 106.200 ;
        RECT 125.400 106.800 125.800 107.200 ;
        RECT 134.200 108.800 134.600 109.200 ;
        RECT 131.000 106.800 131.400 107.200 ;
        RECT 119.000 105.800 119.400 106.200 ;
        RECT 110.200 102.800 110.600 103.200 ;
        RECT 116.600 104.800 117.000 105.200 ;
        RECT 128.600 105.800 129.000 106.200 ;
        RECT 135.000 106.800 135.400 107.200 ;
        RECT 139.800 107.400 140.200 107.800 ;
        RECT 141.400 106.800 141.800 107.200 ;
        RECT 150.200 108.800 150.600 109.200 ;
        RECT 149.400 106.800 149.800 107.200 ;
        RECT 112.600 101.800 113.000 102.200 ;
        RECT 119.000 102.800 119.400 103.200 ;
        RECT 126.200 104.800 126.600 105.200 ;
        RECT 135.800 105.800 136.200 106.200 ;
        RECT 143.800 105.800 144.200 106.200 ;
        RECT 147.000 105.800 147.400 106.200 ;
        RECT 128.600 101.800 129.000 102.200 ;
        RECT 144.600 104.800 145.000 105.200 ;
        RECT 147.000 101.800 147.400 102.200 ;
        RECT 3.000 93.800 3.400 94.200 ;
        RECT 12.600 95.900 13.000 96.300 ;
        RECT 26.200 96.800 26.600 97.200 ;
        RECT 35.800 98.800 36.200 99.200 ;
        RECT 7.000 92.800 7.400 93.200 ;
        RECT 7.800 91.800 8.200 92.200 ;
        RECT 12.600 93.100 13.000 93.500 ;
        RECT 11.000 91.800 11.400 92.200 ;
        RECT 16.600 93.800 17.000 94.200 ;
        RECT 15.000 93.200 15.400 93.600 ;
        RECT 17.400 93.100 17.800 93.500 ;
        RECT 30.200 94.800 30.600 95.200 ;
        RECT 27.800 93.800 28.200 94.200 ;
        RECT 27.000 93.100 27.400 93.500 ;
        RECT 36.600 92.800 37.000 93.200 ;
        RECT 54.200 98.800 54.600 99.200 ;
        RECT 41.400 93.100 41.800 93.500 ;
        RECT 37.400 91.800 37.800 92.200 ;
        RECT 59.800 95.800 60.200 96.200 ;
        RECT 67.800 98.800 68.200 99.200 ;
        RECT 79.000 96.800 79.400 97.200 ;
        RECT 52.600 92.800 53.000 93.200 ;
        RECT 50.200 91.800 50.600 92.200 ;
        RECT 55.800 92.800 56.200 93.200 ;
        RECT 66.200 94.800 66.600 95.200 ;
        RECT 67.800 94.800 68.200 95.200 ;
        RECT 70.200 94.800 70.600 95.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 75.800 95.800 76.200 96.200 ;
        RECT 84.600 98.800 85.000 99.200 ;
        RECT 63.000 92.800 63.400 93.200 ;
        RECT 57.400 91.800 57.800 92.200 ;
        RECT 71.800 91.800 72.200 92.200 ;
        RECT 79.800 94.800 80.200 95.200 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 80.600 93.800 81.000 94.200 ;
        RECT 76.600 92.800 77.000 93.200 ;
        RECT 83.800 93.800 84.200 94.200 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 86.200 93.800 86.600 94.200 ;
        RECT 89.400 98.800 89.800 99.200 ;
        RECT 91.800 98.800 92.200 99.200 ;
        RECT 92.600 96.800 93.000 97.200 ;
        RECT 90.200 93.800 90.600 94.200 ;
        RECT 94.200 93.800 94.600 94.200 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 99.000 95.800 99.400 96.200 ;
        RECT 111.800 98.800 112.200 99.200 ;
        RECT 101.400 94.800 101.800 95.200 ;
        RECT 103.000 94.800 103.400 95.200 ;
        RECT 106.200 92.800 106.600 93.200 ;
        RECT 112.600 96.800 113.000 97.200 ;
        RECT 111.000 95.800 111.400 96.200 ;
        RECT 127.800 98.800 128.200 99.200 ;
        RECT 127.000 96.800 127.400 97.200 ;
        RECT 130.200 96.800 130.600 97.200 ;
        RECT 133.400 96.800 133.800 97.200 ;
        RECT 137.400 96.800 137.800 97.200 ;
        RECT 140.600 96.800 141.000 97.200 ;
        RECT 123.000 95.800 123.400 96.200 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 128.600 95.800 129.000 96.200 ;
        RECT 127.800 94.800 128.200 95.200 ;
        RECT 131.800 95.800 132.200 96.200 ;
        RECT 131.000 94.800 131.400 95.200 ;
        RECT 139.000 95.800 139.400 96.200 ;
        RECT 134.200 94.800 134.600 95.200 ;
        RECT 119.000 92.800 119.400 93.200 ;
        RECT 130.200 91.800 130.600 92.200 ;
        RECT 145.400 93.800 145.800 94.200 ;
        RECT 148.600 96.800 149.000 97.200 ;
        RECT 150.200 95.800 150.600 96.200 ;
        RECT 149.400 94.800 149.800 95.200 ;
        RECT 141.400 91.800 141.800 92.200 ;
        RECT 143.800 91.800 144.200 92.200 ;
        RECT 10.200 88.800 10.600 89.200 ;
        RECT 3.800 84.800 4.200 85.200 ;
        RECT 3.000 83.800 3.400 84.200 ;
        RECT 16.600 88.800 17.000 89.200 ;
        RECT 15.000 87.800 15.400 88.200 ;
        RECT 12.600 81.800 13.000 82.200 ;
        RECT 17.400 86.800 17.800 87.200 ;
        RECT 18.200 85.800 18.600 86.200 ;
        RECT 26.200 87.400 26.600 87.800 ;
        RECT 37.400 88.800 37.800 89.200 ;
        RECT 27.800 86.800 28.200 87.200 ;
        RECT 31.000 85.900 31.400 86.300 ;
        RECT 28.600 85.100 29.000 85.500 ;
        RECT 50.200 86.800 50.600 87.200 ;
        RECT 47.800 85.800 48.200 86.200 ;
        RECT 51.800 85.900 52.200 86.300 ;
        RECT 38.200 85.100 38.600 85.500 ;
        RECT 49.400 85.100 49.800 85.500 ;
        RECT 58.200 81.800 58.600 82.200 ;
        RECT 63.000 88.800 63.400 89.200 ;
        RECT 65.400 88.800 65.800 89.200 ;
        RECT 72.600 88.800 73.000 89.200 ;
        RECT 76.600 88.800 77.000 89.200 ;
        RECT 80.600 88.800 81.000 89.200 ;
        RECT 66.200 84.800 66.600 85.200 ;
        RECT 67.800 84.800 68.200 85.200 ;
        RECT 68.600 84.800 69.000 85.200 ;
        RECT 73.400 86.800 73.800 87.200 ;
        RECT 71.000 85.800 71.400 86.200 ;
        RECT 74.200 85.800 74.600 86.200 ;
        RECT 76.600 84.800 77.000 85.200 ;
        RECT 81.400 86.800 81.800 87.200 ;
        RECT 86.200 88.800 86.600 89.200 ;
        RECT 79.000 84.800 79.400 85.200 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 95.000 86.800 95.400 87.200 ;
        RECT 89.400 84.800 89.800 85.200 ;
        RECT 88.600 82.800 89.000 83.200 ;
        RECT 97.400 86.800 97.800 87.200 ;
        RECT 95.000 85.800 95.400 86.200 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 94.200 84.800 94.600 85.200 ;
        RECT 95.800 81.800 96.200 82.200 ;
        RECT 100.600 84.800 101.000 85.200 ;
        RECT 99.800 81.800 100.200 82.200 ;
        RECT 109.400 86.800 109.800 87.200 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 107.000 84.800 107.400 85.200 ;
        RECT 107.800 81.800 108.200 82.200 ;
        RECT 115.800 86.800 116.200 87.200 ;
        RECT 131.800 88.800 132.200 89.200 ;
        RECT 121.400 86.800 121.800 87.200 ;
        RECT 123.800 85.800 124.200 86.200 ;
        RECT 112.600 81.800 113.000 82.200 ;
        RECT 132.600 86.800 133.000 87.200 ;
        RECT 142.200 88.800 142.600 89.200 ;
        RECT 141.400 86.800 141.800 87.200 ;
        RECT 123.800 83.800 124.200 84.200 ;
        RECT 130.200 84.800 130.600 85.200 ;
        RECT 133.400 85.800 133.800 86.200 ;
        RECT 135.800 85.800 136.200 86.200 ;
        RECT 126.200 81.800 126.600 82.200 ;
        RECT 139.000 85.800 139.400 86.200 ;
        RECT 135.800 81.800 136.200 82.200 ;
        RECT 139.000 81.800 139.400 82.200 ;
        RECT 143.000 81.800 143.400 82.200 ;
        RECT 144.600 81.800 145.000 82.200 ;
        RECT 147.800 81.800 148.200 82.200 ;
        RECT 1.400 71.800 1.800 72.200 ;
        RECT 6.900 75.900 7.300 76.300 ;
        RECT 3.800 72.800 4.200 73.200 ;
        RECT 4.600 71.800 5.000 72.200 ;
        RECT 6.900 73.100 7.300 73.500 ;
        RECT 28.600 75.800 29.000 76.200 ;
        RECT 15.000 74.800 15.400 75.200 ;
        RECT 9.400 71.800 9.800 72.200 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 17.400 71.800 17.800 72.200 ;
        RECT 19.800 73.100 20.200 73.500 ;
        RECT 59.000 76.800 59.400 77.200 ;
        RECT 29.400 73.100 29.800 73.500 ;
        RECT 38.200 73.800 38.600 74.200 ;
        RECT 39.000 73.100 39.400 73.500 ;
        RECT 47.800 71.800 48.200 72.200 ;
        RECT 50.200 73.100 50.600 73.500 ;
        RECT 59.800 73.800 60.200 74.200 ;
        RECT 52.600 72.800 53.000 73.200 ;
        RECT 64.600 76.800 65.000 77.200 ;
        RECT 64.600 75.800 65.000 76.200 ;
        RECT 63.800 74.800 64.200 75.200 ;
        RECT 75.800 78.800 76.200 79.200 ;
        RECT 71.000 72.800 71.400 73.200 ;
        RECT 66.200 71.800 66.600 72.200 ;
        RECT 79.800 73.800 80.200 74.200 ;
        RECT 75.800 71.800 76.200 72.200 ;
        RECT 83.800 73.800 84.200 74.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 91.800 72.800 92.200 73.200 ;
        RECT 97.400 73.800 97.800 74.200 ;
        RECT 85.400 71.800 85.800 72.200 ;
        RECT 87.800 71.800 88.200 72.200 ;
        RECT 94.200 71.800 94.600 72.200 ;
        RECT 106.200 76.800 106.600 77.200 ;
        RECT 98.200 71.800 98.600 72.200 ;
        RECT 103.000 71.800 103.400 72.200 ;
        RECT 107.000 72.800 107.400 73.200 ;
        RECT 109.400 73.800 109.800 74.200 ;
        RECT 118.200 78.800 118.600 79.200 ;
        RECT 112.600 76.800 113.000 77.200 ;
        RECT 115.800 76.800 116.200 77.200 ;
        RECT 114.200 75.800 114.600 76.200 ;
        RECT 113.400 74.800 113.800 75.200 ;
        RECT 121.400 76.800 121.800 77.200 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 107.800 71.800 108.200 72.200 ;
        RECT 111.000 71.800 111.400 72.200 ;
        RECT 115.800 71.800 116.200 72.200 ;
        RECT 119.800 75.800 120.200 76.200 ;
        RECT 127.800 76.800 128.200 77.200 ;
        RECT 126.200 75.800 126.600 76.200 ;
        RECT 119.000 73.800 119.400 74.200 ;
        RECT 130.200 74.800 130.600 75.200 ;
        RECT 133.300 75.900 133.700 76.300 ;
        RECT 139.800 76.800 140.200 77.200 ;
        RECT 145.400 76.800 145.800 77.200 ;
        RECT 141.400 75.800 141.800 76.200 ;
        RECT 125.400 73.800 125.800 74.200 ;
        RECT 133.300 73.100 133.700 73.500 ;
        RECT 137.400 73.800 137.800 74.200 ;
        RECT 147.000 75.800 147.400 76.200 ;
        RECT 150.200 78.800 150.600 79.200 ;
        RECT 146.200 74.800 146.600 75.200 ;
        RECT 143.800 71.800 144.200 72.200 ;
        RECT 145.400 71.800 145.800 72.200 ;
        RECT 11.000 66.800 11.400 67.200 ;
        RECT 13.400 65.800 13.800 66.200 ;
        RECT 5.400 61.800 5.800 62.200 ;
        RECT 12.600 61.800 13.000 62.200 ;
        RECT 15.800 64.800 16.200 65.200 ;
        RECT 21.400 68.800 21.800 69.200 ;
        RECT 21.400 67.400 21.800 67.800 ;
        RECT 27.000 68.800 27.400 69.200 ;
        RECT 23.000 66.800 23.400 67.200 ;
        RECT 27.000 67.400 27.400 67.800 ;
        RECT 28.600 66.800 29.000 67.200 ;
        RECT 32.600 67.400 33.000 67.800 ;
        RECT 57.400 68.800 57.800 69.200 ;
        RECT 36.600 65.800 37.000 66.200 ;
        RECT 39.800 65.900 40.200 66.300 ;
        RECT 37.400 65.100 37.800 65.500 ;
        RECT 49.400 66.800 49.800 67.200 ;
        RECT 59.800 68.800 60.200 69.200 ;
        RECT 52.600 66.800 53.000 67.200 ;
        RECT 51.000 65.900 51.400 66.300 ;
        RECT 46.200 61.800 46.600 62.200 ;
        RECT 48.600 65.100 49.000 65.500 ;
        RECT 67.800 67.800 68.200 68.200 ;
        RECT 60.600 64.800 61.000 65.200 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 62.200 64.800 62.600 65.200 ;
        RECT 67.800 65.800 68.200 66.200 ;
        RECT 77.400 65.800 77.800 66.200 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 64.600 62.800 65.000 63.200 ;
        RECT 76.600 64.800 77.000 65.200 ;
        RECT 79.000 64.800 79.400 65.200 ;
        RECT 87.000 68.800 87.400 69.200 ;
        RECT 81.400 64.800 81.800 65.200 ;
        RECT 85.400 65.800 85.800 66.200 ;
        RECT 88.600 64.800 89.000 65.200 ;
        RECT 94.200 66.800 94.600 67.200 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 97.400 65.800 97.800 66.200 ;
        RECT 112.600 68.800 113.000 69.200 ;
        RECT 107.800 66.800 108.200 67.200 ;
        RECT 104.600 65.800 105.000 66.200 ;
        RECT 110.200 64.800 110.600 65.200 ;
        RECT 106.200 61.800 106.600 62.200 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 115.000 61.800 115.400 62.200 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 124.600 66.800 125.000 67.200 ;
        RECT 138.200 68.800 138.600 69.200 ;
        RECT 117.400 61.800 117.800 62.200 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 149.400 67.400 149.800 67.800 ;
        RECT 141.400 65.800 141.800 66.200 ;
        RECT 131.000 61.800 131.400 62.200 ;
        RECT 134.200 61.800 134.600 62.200 ;
        RECT 151.000 66.800 151.400 67.200 ;
        RECT 144.600 65.800 145.000 66.200 ;
        RECT 139.800 61.800 140.200 62.200 ;
        RECT 143.000 61.800 143.400 62.200 ;
        RECT 149.400 61.800 149.800 62.200 ;
        RECT 1.300 55.900 1.700 56.300 ;
        RECT 19.000 58.800 19.400 59.200 ;
        RECT 16.500 55.900 16.900 56.300 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 1.300 53.100 1.700 53.500 ;
        RECT 5.400 53.800 5.800 54.200 ;
        RECT 6.200 53.100 6.600 53.500 ;
        RECT 15.000 51.800 15.400 52.200 ;
        RECT 16.500 53.100 16.900 53.500 ;
        RECT 20.600 53.800 21.000 54.200 ;
        RECT 21.400 53.800 21.800 54.200 ;
        RECT 23.800 55.800 24.200 56.200 ;
        RECT 24.600 55.800 25.000 56.200 ;
        RECT 31.000 58.800 31.400 59.200 ;
        RECT 25.400 52.800 25.800 53.200 ;
        RECT 47.800 58.800 48.200 59.200 ;
        RECT 42.200 54.800 42.600 55.200 ;
        RECT 52.600 58.800 53.000 59.200 ;
        RECT 55.000 58.800 55.400 59.200 ;
        RECT 39.800 53.800 40.200 54.200 ;
        RECT 39.000 53.100 39.400 53.500 ;
        RECT 55.000 55.800 55.400 56.200 ;
        RECT 55.800 55.800 56.200 56.200 ;
        RECT 51.000 53.800 51.400 54.200 ;
        RECT 55.000 54.800 55.400 55.200 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 61.400 53.800 61.800 54.200 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 68.600 53.800 69.000 54.200 ;
        RECT 58.200 51.800 58.600 52.200 ;
        RECT 60.600 51.800 61.000 52.200 ;
        RECT 63.000 51.800 63.400 52.200 ;
        RECT 64.600 51.800 65.000 52.200 ;
        RECT 72.600 53.800 73.000 54.200 ;
        RECT 74.200 53.800 74.600 54.200 ;
        RECT 76.600 53.800 77.000 54.200 ;
        RECT 77.400 53.800 77.800 54.200 ;
        RECT 79.800 56.800 80.200 57.200 ;
        RECT 93.400 56.800 93.800 57.200 ;
        RECT 95.800 56.800 96.200 57.200 ;
        RECT 91.800 55.800 92.200 56.200 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 82.200 53.800 82.600 54.200 ;
        RECT 80.600 52.800 81.000 53.200 ;
        RECT 82.200 52.800 82.600 53.200 ;
        RECT 75.800 51.800 76.200 52.200 ;
        RECT 79.000 51.800 79.400 52.200 ;
        RECT 83.000 51.800 83.400 52.200 ;
        RECT 87.000 52.800 87.400 53.200 ;
        RECT 97.400 55.800 97.800 56.200 ;
        RECT 107.000 56.800 107.400 57.200 ;
        RECT 96.600 54.800 97.000 55.200 ;
        RECT 89.400 51.800 89.800 52.200 ;
        RECT 108.600 55.800 109.000 56.200 ;
        RECT 114.200 56.800 114.600 57.200 ;
        RECT 116.600 56.800 117.000 57.200 ;
        RECT 107.800 54.800 108.200 55.200 ;
        RECT 112.600 55.800 113.000 56.200 ;
        RECT 96.600 51.800 97.000 52.200 ;
        RECT 99.800 51.800 100.200 52.200 ;
        RECT 118.200 55.800 118.600 56.200 ;
        RECT 123.000 56.800 123.400 57.200 ;
        RECT 117.400 54.800 117.800 55.200 ;
        RECT 111.000 51.800 111.400 52.200 ;
        RECT 115.000 51.800 115.400 52.200 ;
        RECT 124.600 55.800 125.000 56.200 ;
        RECT 136.600 56.800 137.000 57.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 120.600 51.800 121.000 52.200 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 135.000 55.800 135.400 56.200 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 126.200 52.800 126.600 53.200 ;
        RECT 138.200 53.800 138.600 54.200 ;
        RECT 137.400 51.800 137.800 52.200 ;
        RECT 143.000 55.900 143.400 56.300 ;
        RECT 140.600 51.800 141.000 52.200 ;
        RECT 143.000 53.100 143.400 53.500 ;
        RECT 148.600 54.800 149.000 55.200 ;
        RECT 147.000 53.800 147.400 54.200 ;
        RECT 145.400 53.200 145.800 53.600 ;
        RECT 145.400 51.800 145.800 52.200 ;
        RECT 8.600 48.800 9.000 49.200 ;
        RECT 15.000 47.400 15.400 47.800 ;
        RECT 26.200 48.800 26.600 49.200 ;
        RECT 3.000 45.800 3.400 46.200 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 18.200 46.800 18.600 47.200 ;
        RECT 19.800 45.900 20.200 46.300 ;
        RECT 17.400 45.100 17.800 45.500 ;
        RECT 6.200 43.800 6.600 44.200 ;
        RECT 34.200 45.800 34.600 46.200 ;
        RECT 43.000 47.800 43.400 48.200 ;
        RECT 39.800 45.800 40.200 46.200 ;
        RECT 42.200 44.800 42.600 45.200 ;
        RECT 47.800 48.800 48.200 49.200 ;
        RECT 44.600 46.800 45.000 47.200 ;
        RECT 47.000 46.800 47.400 47.200 ;
        RECT 46.200 45.800 46.600 46.200 ;
        RECT 48.600 46.800 49.000 47.200 ;
        RECT 55.000 47.400 55.400 47.800 ;
        RECT 66.200 48.800 66.600 49.200 ;
        RECT 56.600 46.800 57.000 47.200 ;
        RECT 49.400 45.800 49.800 46.200 ;
        RECT 59.800 45.900 60.200 46.300 ;
        RECT 57.400 45.100 57.800 45.500 ;
        RECT 81.400 48.800 81.800 49.200 ;
        RECT 88.600 47.800 89.000 48.200 ;
        RECT 92.600 48.800 93.000 49.200 ;
        RECT 78.200 44.800 78.600 45.200 ;
        RECT 75.800 43.800 76.200 44.200 ;
        RECT 87.800 45.800 88.200 46.200 ;
        RECT 90.200 45.800 90.600 46.200 ;
        RECT 103.800 48.800 104.200 49.200 ;
        RECT 105.400 45.800 105.800 46.200 ;
        RECT 92.600 41.800 93.000 42.200 ;
        RECT 99.800 41.800 100.200 42.200 ;
        RECT 116.600 48.800 117.000 49.200 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 115.000 45.800 115.400 46.200 ;
        RECT 117.400 46.800 117.800 47.200 ;
        RECT 123.000 48.800 123.400 49.200 ;
        RECT 110.200 44.800 110.600 45.200 ;
        RECT 114.200 44.800 114.600 45.200 ;
        RECT 118.200 45.800 118.600 46.200 ;
        RECT 119.800 41.800 120.200 42.200 ;
        RECT 124.600 46.800 125.000 47.200 ;
        RECT 134.200 48.800 134.600 49.200 ;
        RECT 128.600 45.800 129.000 46.200 ;
        RECT 131.800 45.800 132.200 46.200 ;
        RECT 135.000 46.800 135.400 47.200 ;
        RECT 126.200 41.800 126.600 42.200 ;
        RECT 129.400 44.800 129.800 45.200 ;
        RECT 135.800 45.800 136.200 46.200 ;
        RECT 130.200 41.800 130.600 42.200 ;
        RECT 131.800 41.800 132.200 42.200 ;
        RECT 141.400 44.800 141.800 45.200 ;
        RECT 143.000 41.800 143.400 42.200 ;
        RECT 147.800 43.800 148.200 44.200 ;
        RECT 150.200 41.800 150.600 42.200 ;
        RECT 1.500 35.900 1.900 36.300 ;
        RECT 2.100 34.900 2.500 35.300 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 14.200 35.900 14.600 36.300 ;
        RECT 3.800 34.800 4.200 35.200 ;
        RECT 1.500 33.100 1.900 33.500 ;
        RECT 16.600 35.800 17.000 36.200 ;
        RECT 27.800 38.800 28.200 39.200 ;
        RECT 12.600 33.800 13.000 34.200 ;
        RECT 14.200 33.100 14.600 33.500 ;
        RECT 10.200 31.800 10.600 32.200 ;
        RECT 18.200 33.800 18.600 34.200 ;
        RECT 16.600 33.200 17.000 33.600 ;
        RECT 19.000 33.100 19.400 33.500 ;
        RECT 37.400 34.800 37.800 35.200 ;
        RECT 21.400 32.800 21.800 33.200 ;
        RECT 28.600 33.100 29.000 33.500 ;
        RECT 31.000 32.800 31.400 33.200 ;
        RECT 38.200 38.800 38.600 39.200 ;
        RECT 40.600 35.900 41.000 36.300 ;
        RECT 43.000 35.800 43.400 36.200 ;
        RECT 46.200 38.800 46.600 39.200 ;
        RECT 39.800 33.800 40.200 34.200 ;
        RECT 40.600 33.100 41.000 33.500 ;
        RECT 44.600 33.800 45.000 34.200 ;
        RECT 43.000 33.200 43.400 33.600 ;
        RECT 52.600 38.800 53.000 39.200 ;
        RECT 50.300 35.900 50.700 36.300 ;
        RECT 63.800 38.800 64.200 39.200 ;
        RECT 50.900 34.900 51.300 35.300 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 58.200 34.800 58.600 35.200 ;
        RECT 50.300 33.100 50.700 33.500 ;
        RECT 54.200 33.800 54.600 34.200 ;
        RECT 55.000 33.100 55.400 33.500 ;
        RECT 57.400 32.800 57.800 33.200 ;
        RECT 65.400 33.800 65.800 34.200 ;
        RECT 64.600 33.100 65.000 33.500 ;
        RECT 79.800 38.800 80.200 39.200 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 74.200 33.800 74.600 34.200 ;
        RECT 73.400 31.800 73.800 32.200 ;
        RECT 78.200 32.800 78.600 33.200 ;
        RECT 79.000 32.800 79.400 33.200 ;
        RECT 81.400 34.800 81.800 35.200 ;
        RECT 87.800 34.800 88.200 35.200 ;
        RECT 91.000 34.800 91.400 35.200 ;
        RECT 83.000 31.800 83.400 32.200 ;
        RECT 85.400 32.800 85.800 33.200 ;
        RECT 88.600 33.800 89.000 34.200 ;
        RECT 84.600 31.800 85.000 32.200 ;
        RECT 86.200 31.800 86.600 32.200 ;
        RECT 89.400 32.800 89.800 33.200 ;
        RECT 93.400 32.800 93.800 33.200 ;
        RECT 111.000 36.800 111.400 37.200 ;
        RECT 109.400 35.800 109.800 36.200 ;
        RECT 103.800 33.800 104.200 34.200 ;
        RECT 95.800 31.800 96.200 32.200 ;
        RECT 104.600 32.800 105.000 33.200 ;
        RECT 112.600 34.800 113.000 35.200 ;
        RECT 113.400 34.800 113.800 35.200 ;
        RECT 107.000 32.800 107.400 33.200 ;
        RECT 119.000 34.800 119.400 35.200 ;
        RECT 118.200 33.800 118.600 34.200 ;
        RECT 122.200 34.800 122.600 35.200 ;
        RECT 130.200 35.800 130.600 36.200 ;
        RECT 131.000 35.800 131.400 36.200 ;
        RECT 138.200 36.800 138.600 37.200 ;
        RECT 145.400 36.800 145.800 37.200 ;
        RECT 120.600 33.800 121.000 34.200 ;
        RECT 124.600 33.800 125.000 34.200 ;
        RECT 116.600 31.800 117.000 32.200 ;
        RECT 125.400 31.800 125.800 32.200 ;
        RECT 139.000 34.800 139.400 35.200 ;
        RECT 143.800 35.800 144.200 36.200 ;
        RECT 148.600 34.800 149.000 35.200 ;
        RECT 150.200 33.800 150.600 34.200 ;
        RECT 147.000 31.800 147.400 32.200 ;
        RECT 11.000 27.400 11.400 27.800 ;
        RECT 22.200 28.800 22.600 29.200 ;
        RECT 14.200 26.800 14.600 27.200 ;
        RECT 31.800 28.800 32.200 29.200 ;
        RECT 15.800 25.900 16.200 26.300 ;
        RECT 13.400 25.100 13.800 25.500 ;
        RECT 6.200 21.800 6.600 22.200 ;
        RECT 23.800 26.800 24.200 27.200 ;
        RECT 41.400 28.800 41.800 29.200 ;
        RECT 25.400 25.900 25.800 26.300 ;
        RECT 20.600 23.800 21.000 24.200 ;
        RECT 23.000 25.100 23.400 25.500 ;
        RECT 33.400 26.800 33.800 27.200 ;
        RECT 51.000 28.800 51.400 29.200 ;
        RECT 35.000 25.900 35.400 26.300 ;
        RECT 32.600 25.100 33.000 25.500 ;
        RECT 62.200 28.800 62.600 29.200 ;
        RECT 44.600 25.900 45.000 26.300 ;
        RECT 42.200 25.100 42.600 25.500 ;
        RECT 57.400 26.800 57.800 27.200 ;
        RECT 55.800 25.900 56.200 26.300 ;
        RECT 53.400 25.100 53.800 25.500 ;
        RECT 79.000 27.400 79.400 27.800 ;
        RECT 63.800 21.800 64.200 22.200 ;
        RECT 75.800 21.800 76.200 22.200 ;
        RECT 79.800 21.800 80.200 22.200 ;
        RECT 91.000 28.800 91.400 29.200 ;
        RECT 86.200 26.800 86.600 27.200 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 87.000 25.800 87.400 26.200 ;
        RECT 87.800 25.800 88.200 26.200 ;
        RECT 97.400 26.800 97.800 27.200 ;
        RECT 103.800 28.800 104.200 29.200 ;
        RECT 97.400 25.800 97.800 26.200 ;
        RECT 99.800 25.800 100.200 26.200 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 105.400 25.800 105.800 26.200 ;
        RECT 107.800 25.800 108.200 26.200 ;
        RECT 108.600 25.800 109.000 26.200 ;
        RECT 99.800 22.800 100.200 23.200 ;
        RECT 112.600 25.800 113.000 26.200 ;
        RECT 121.400 27.800 121.800 28.200 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 119.000 26.800 119.400 27.200 ;
        RECT 120.600 26.800 121.000 27.200 ;
        RECT 106.200 21.800 106.600 22.200 ;
        RECT 123.000 25.800 123.400 26.200 ;
        RECT 126.200 25.800 126.600 26.200 ;
        RECT 115.800 21.800 116.200 22.200 ;
        RECT 125.400 24.800 125.800 25.200 ;
        RECT 129.400 26.800 129.800 27.200 ;
        RECT 127.800 25.800 128.200 26.200 ;
        RECT 131.800 25.800 132.200 26.200 ;
        RECT 132.600 25.800 133.000 26.200 ;
        RECT 134.200 25.800 134.600 26.200 ;
        RECT 131.000 24.800 131.400 25.200 ;
        RECT 136.600 25.800 137.000 26.200 ;
        RECT 139.800 25.800 140.200 26.200 ;
        RECT 140.600 24.800 141.000 25.200 ;
        RECT 141.400 24.800 141.800 25.200 ;
        RECT 147.000 28.800 147.400 29.200 ;
        RECT 142.200 21.800 142.600 22.200 ;
        RECT 144.600 22.800 145.000 23.200 ;
        RECT 9.400 18.800 9.800 19.200 ;
        RECT 0.600 13.100 1.000 13.500 ;
        RECT 12.500 15.900 12.900 16.300 ;
        RECT 26.200 18.800 26.600 19.200 ;
        RECT 11.000 11.800 11.400 12.200 ;
        RECT 12.500 13.100 12.900 13.500 ;
        RECT 30.200 18.800 30.600 19.200 ;
        RECT 27.700 15.900 28.100 16.300 ;
        RECT 41.400 16.800 41.800 17.200 ;
        RECT 17.400 13.100 17.800 13.500 ;
        RECT 36.600 14.800 37.000 15.200 ;
        RECT 27.700 13.100 28.100 13.500 ;
        RECT 31.800 13.800 32.200 14.200 ;
        RECT 33.400 13.800 33.800 14.200 ;
        RECT 32.600 13.100 33.000 13.500 ;
        RECT 60.600 16.800 61.000 17.200 ;
        RECT 70.200 18.800 70.600 19.200 ;
        RECT 45.400 13.800 45.800 14.200 ;
        RECT 47.000 12.800 47.400 13.200 ;
        RECT 51.800 13.100 52.200 13.500 ;
        RECT 64.600 14.800 65.000 15.200 ;
        RECT 54.200 12.800 54.600 13.200 ;
        RECT 61.400 13.100 61.800 13.500 ;
        RECT 72.600 16.800 73.000 17.200 ;
        RECT 71.000 13.800 71.400 14.200 ;
        RECT 76.600 15.800 77.000 16.200 ;
        RECT 75.000 12.800 75.400 13.200 ;
        RECT 78.200 14.800 78.600 15.200 ;
        RECT 79.800 11.800 80.200 12.200 ;
        RECT 82.200 12.800 82.600 13.200 ;
        RECT 87.800 14.000 88.200 14.400 ;
        RECT 95.800 16.800 96.200 17.200 ;
        RECT 94.200 15.800 94.600 16.200 ;
        RECT 104.600 18.800 105.000 19.200 ;
        RECT 103.800 16.800 104.200 17.200 ;
        RECT 91.800 12.800 92.200 13.200 ;
        RECT 97.400 12.800 97.800 13.200 ;
        RECT 98.200 11.800 98.600 12.200 ;
        RECT 105.400 15.800 105.800 16.200 ;
        RECT 109.400 16.800 109.800 17.200 ;
        RECT 104.600 14.800 105.000 15.200 ;
        RECT 106.200 14.800 106.600 15.200 ;
        RECT 102.200 12.800 102.600 13.200 ;
        RECT 109.400 14.800 109.800 15.200 ;
        RECT 107.000 12.800 107.400 13.200 ;
        RECT 110.200 13.800 110.600 14.200 ;
        RECT 128.600 18.800 129.000 19.200 ;
        RECT 132.600 16.800 133.000 17.200 ;
        RECT 126.200 15.800 126.600 16.200 ;
        RECT 130.200 15.900 130.600 16.300 ;
        RECT 120.600 12.800 121.000 13.200 ;
        RECT 121.400 12.800 121.800 13.200 ;
        RECT 113.400 11.800 113.800 12.200 ;
        RECT 123.800 12.800 124.200 13.200 ;
        RECT 124.600 11.800 125.000 12.200 ;
        RECT 130.200 13.100 130.600 13.500 ;
        RECT 134.200 13.800 134.600 14.200 ;
        RECT 135.800 13.800 136.200 14.200 ;
        RECT 132.600 13.200 133.000 13.600 ;
        RECT 135.000 13.100 135.400 13.500 ;
        RECT 3.800 8.800 4.200 9.200 ;
        RECT 8.600 8.800 9.000 9.200 ;
        RECT 15.000 8.800 15.400 9.200 ;
        RECT 15.000 7.400 15.400 7.800 ;
        RECT 7.800 4.800 8.200 5.200 ;
        RECT 16.600 6.800 17.000 7.200 ;
        RECT 25.400 8.800 25.800 9.200 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 51.000 8.800 51.400 9.200 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 44.600 6.800 45.000 7.200 ;
        RECT 40.600 5.100 41.000 5.500 ;
        RECT 51.800 5.100 52.200 5.500 ;
        RECT 71.800 6.800 72.200 7.200 ;
        RECT 66.200 6.100 66.600 6.500 ;
        RECT 70.200 5.900 70.600 6.300 ;
        RECT 80.600 6.800 81.000 7.200 ;
        RECT 78.200 6.100 78.600 6.500 ;
        RECT 72.600 5.100 73.000 5.500 ;
        RECT 82.200 5.900 82.600 6.300 ;
        RECT 87.800 5.900 88.200 6.300 ;
        RECT 84.600 5.100 85.000 5.500 ;
        RECT 85.400 5.100 85.800 5.500 ;
        RECT 99.800 6.800 100.200 7.200 ;
        RECT 101.400 5.900 101.800 6.300 ;
        RECT 99.000 5.100 99.400 5.500 ;
        RECT 111.800 6.800 112.200 7.200 ;
        RECT 113.400 5.900 113.800 6.300 ;
        RECT 111.000 5.100 111.400 5.500 ;
        RECT 123.800 6.800 124.200 7.200 ;
        RECT 125.400 5.900 125.800 6.300 ;
        RECT 123.000 5.100 123.400 5.500 ;
        RECT 135.800 6.800 136.200 7.200 ;
        RECT 135.000 5.100 135.400 5.500 ;
        RECT 147.000 4.800 147.400 5.200 ;
      LAYER metal2 ;
        RECT 17.400 128.800 17.800 129.200 ;
        RECT 29.400 129.100 29.800 129.200 ;
        RECT 30.200 129.100 30.600 129.200 ;
        RECT 29.400 128.800 30.600 129.100 ;
        RECT 0.600 128.100 1.000 128.200 ;
        RECT 1.400 128.100 1.800 128.200 ;
        RECT 0.600 127.800 1.800 128.100 ;
        RECT 5.400 128.100 5.800 128.200 ;
        RECT 6.200 128.100 6.600 128.200 ;
        RECT 5.400 127.800 6.600 128.100 ;
        RECT 7.800 127.800 8.200 128.200 ;
        RECT 6.200 126.800 6.600 127.200 ;
        RECT 6.200 126.200 6.500 126.800 ;
        RECT 7.800 126.200 8.100 127.800 ;
        RECT 12.600 127.500 13.000 127.900 ;
        RECT 15.700 127.800 16.100 127.900 ;
        RECT 13.300 127.500 16.100 127.800 ;
        RECT 8.600 126.800 9.000 127.200 ;
        RECT 10.200 127.100 10.600 127.200 ;
        RECT 11.000 127.100 11.400 127.200 ;
        RECT 10.200 126.800 11.400 127.100 ;
        RECT 12.600 127.100 12.900 127.500 ;
        RECT 13.300 127.400 13.700 127.500 ;
        RECT 15.000 127.400 15.400 127.500 ;
        RECT 12.600 126.800 15.400 127.100 ;
        RECT 8.600 126.200 8.900 126.800 ;
        RECT 6.200 125.800 6.600 126.200 ;
        RECT 7.000 126.100 7.400 126.200 ;
        RECT 7.800 126.100 8.200 126.200 ;
        RECT 7.000 125.800 8.200 126.100 ;
        RECT 8.600 125.800 9.000 126.200 ;
        RECT 9.400 125.800 9.800 126.200 ;
        RECT 10.200 126.100 10.600 126.200 ;
        RECT 11.000 126.100 11.400 126.200 ;
        RECT 10.200 125.800 11.400 126.100 ;
        RECT 3.800 115.900 4.200 116.300 ;
        RECT 6.900 115.900 7.300 116.300 ;
        RECT 3.800 114.200 4.100 115.900 ;
        RECT 6.300 114.900 6.700 115.300 ;
        RECT 6.300 114.200 6.600 114.900 ;
        RECT 3.800 113.900 6.600 114.200 ;
        RECT 3.800 113.500 4.100 113.900 ;
        RECT 4.500 113.500 4.900 113.600 ;
        RECT 6.200 113.500 6.600 113.600 ;
        RECT 7.000 113.500 7.300 115.900 ;
        RECT 9.400 114.200 9.700 125.800 ;
        RECT 12.600 125.100 12.900 126.800 ;
        RECT 13.400 126.100 13.800 126.200 ;
        RECT 14.200 126.100 14.600 126.200 ;
        RECT 13.400 125.800 14.600 126.100 ;
        RECT 15.100 126.100 15.400 126.800 ;
        RECT 15.100 125.700 15.500 126.100 ;
        RECT 15.800 125.100 16.100 127.500 ;
        RECT 16.600 126.800 17.000 127.200 ;
        RECT 16.600 126.200 16.900 126.800 ;
        RECT 16.600 125.800 17.000 126.200 ;
        RECT 12.600 124.700 13.000 125.100 ;
        RECT 15.700 124.700 16.100 125.100 ;
        RECT 17.400 125.200 17.700 128.800 ;
        RECT 24.600 127.500 25.000 127.900 ;
        RECT 27.700 127.800 28.100 127.900 ;
        RECT 25.300 127.500 28.100 127.800 ;
        RECT 19.800 127.100 20.200 127.200 ;
        RECT 20.600 127.100 21.000 127.200 ;
        RECT 19.800 126.800 21.000 127.100 ;
        RECT 21.400 126.800 21.800 127.200 ;
        RECT 24.600 127.100 24.900 127.500 ;
        RECT 25.300 127.400 25.700 127.500 ;
        RECT 27.000 127.400 27.400 127.500 ;
        RECT 24.600 126.800 27.400 127.100 ;
        RECT 21.400 126.200 21.700 126.800 ;
        RECT 21.400 125.800 21.800 126.200 ;
        RECT 17.400 124.800 17.800 125.200 ;
        RECT 24.600 125.100 24.900 126.800 ;
        RECT 27.100 126.100 27.400 126.800 ;
        RECT 27.100 125.700 27.500 126.100 ;
        RECT 26.200 125.100 26.600 125.200 ;
        RECT 27.000 125.100 27.400 125.200 ;
        RECT 27.800 125.100 28.100 127.500 ;
        RECT 31.000 126.800 31.400 127.200 ;
        RECT 31.000 125.200 31.300 126.800 ;
        RECT 24.600 124.700 25.000 125.100 ;
        RECT 26.200 124.800 27.400 125.100 ;
        RECT 27.700 124.700 28.100 125.100 ;
        RECT 28.600 125.100 29.000 125.200 ;
        RECT 29.400 125.100 29.800 125.200 ;
        RECT 28.600 124.800 29.800 125.100 ;
        RECT 30.200 124.800 30.600 125.200 ;
        RECT 31.000 124.800 31.400 125.200 ;
        RECT 31.800 125.100 32.200 127.900 ;
        RECT 11.800 115.900 12.200 116.300 ;
        RECT 15.100 115.900 15.500 116.300 ;
        RECT 10.200 114.800 10.600 115.200 ;
        RECT 9.400 113.800 9.800 114.200 ;
        RECT 3.800 113.100 4.200 113.500 ;
        RECT 4.500 113.200 7.300 113.500 ;
        RECT 6.900 113.100 7.300 113.200 ;
        RECT 8.600 112.800 9.000 113.200 ;
        RECT 2.200 111.800 2.600 112.200 ;
        RECT 5.400 112.100 5.800 112.200 ;
        RECT 6.200 112.100 6.600 112.200 ;
        RECT 5.400 111.800 6.600 112.100 ;
        RECT 7.000 111.800 7.400 112.200 ;
        RECT 1.400 110.800 1.800 111.200 ;
        RECT 1.400 109.200 1.700 110.800 ;
        RECT 2.200 110.200 2.500 111.800 ;
        RECT 2.200 109.800 2.600 110.200 ;
        RECT 7.000 109.200 7.300 111.800 ;
        RECT 8.600 111.200 8.900 112.800 ;
        RECT 10.200 112.200 10.500 114.800 ;
        RECT 11.800 114.200 12.100 115.900 ;
        RECT 13.800 114.200 14.200 114.300 ;
        RECT 11.800 113.900 14.200 114.200 ;
        RECT 11.800 113.500 12.100 113.900 ;
        RECT 12.500 113.500 12.900 113.600 ;
        RECT 14.200 113.500 14.600 113.600 ;
        RECT 15.200 113.500 15.500 115.900 ;
        RECT 16.600 116.100 17.000 116.200 ;
        RECT 17.400 116.100 17.800 116.200 ;
        RECT 16.600 115.800 17.800 116.100 ;
        RECT 19.800 116.100 20.200 116.200 ;
        RECT 20.600 116.100 21.000 116.200 ;
        RECT 19.800 115.800 21.000 116.100 ;
        RECT 24.600 115.900 25.000 116.300 ;
        RECT 26.200 116.100 26.600 116.200 ;
        RECT 27.000 116.100 27.400 116.200 ;
        RECT 15.800 114.800 16.200 115.200 ;
        RECT 19.000 114.800 19.400 115.200 ;
        RECT 15.800 114.200 16.100 114.800 ;
        RECT 15.800 113.800 16.200 114.200 ;
        RECT 17.400 114.100 17.800 114.200 ;
        RECT 18.200 114.100 18.600 114.200 ;
        RECT 17.400 113.800 18.600 114.100 ;
        RECT 11.800 113.100 12.200 113.500 ;
        RECT 12.500 113.200 14.600 113.500 ;
        RECT 15.100 113.100 15.500 113.500 ;
        RECT 16.600 112.800 17.000 113.200 ;
        RECT 16.600 112.200 16.900 112.800 ;
        RECT 10.200 111.800 10.600 112.200 ;
        RECT 13.400 111.800 13.800 112.200 ;
        RECT 16.600 111.800 17.000 112.200 ;
        RECT 8.600 110.800 9.000 111.200 ;
        RECT 8.600 109.800 9.000 110.200 ;
        RECT 1.400 108.800 1.800 109.200 ;
        RECT 3.800 108.800 4.200 109.200 ;
        RECT 7.000 108.800 7.400 109.200 ;
        RECT 3.800 108.200 4.100 108.800 ;
        RECT 3.800 107.800 4.200 108.200 ;
        RECT 7.000 108.100 7.400 108.200 ;
        RECT 7.800 108.100 8.200 108.200 ;
        RECT 7.000 107.800 8.200 108.100 ;
        RECT 8.600 107.200 8.900 109.800 ;
        RECT 8.600 106.800 9.000 107.200 ;
        RECT 10.200 105.800 10.600 106.200 ;
        RECT 10.200 105.200 10.500 105.800 ;
        RECT 10.200 104.800 10.600 105.200 ;
        RECT 11.000 105.100 11.400 107.900 ;
        RECT 12.600 103.100 13.000 108.900 ;
        RECT 13.400 106.300 13.700 111.800 ;
        RECT 19.000 111.200 19.300 114.800 ;
        RECT 24.600 114.200 24.900 115.900 ;
        RECT 26.200 115.800 27.400 116.100 ;
        RECT 27.700 115.900 28.100 116.300 ;
        RECT 27.100 114.900 27.500 115.300 ;
        RECT 27.100 114.200 27.400 114.900 ;
        RECT 20.600 114.100 21.000 114.200 ;
        RECT 21.400 114.100 21.800 114.200 ;
        RECT 20.600 113.800 21.800 114.100 ;
        RECT 23.000 113.800 23.400 114.200 ;
        RECT 24.600 113.900 27.400 114.200 ;
        RECT 23.000 113.200 23.300 113.800 ;
        RECT 24.600 113.500 24.900 113.900 ;
        RECT 25.300 113.500 25.700 113.600 ;
        RECT 27.000 113.500 27.400 113.600 ;
        RECT 27.800 113.500 28.100 115.900 ;
        RECT 28.600 114.800 29.000 115.200 ;
        RECT 28.600 114.200 28.900 114.800 ;
        RECT 28.600 113.800 29.000 114.200 ;
        RECT 23.000 112.800 23.400 113.200 ;
        RECT 24.600 113.100 25.000 113.500 ;
        RECT 25.300 113.200 28.100 113.500 ;
        RECT 27.700 113.100 28.100 113.200 ;
        RECT 29.400 113.100 29.800 115.900 ;
        RECT 21.400 111.800 21.800 112.200 ;
        RECT 19.000 110.800 19.400 111.200 ;
        RECT 19.800 109.100 20.200 109.200 ;
        RECT 20.600 109.100 21.000 109.200 ;
        RECT 16.600 106.800 17.000 107.200 ;
        RECT 13.400 105.900 13.800 106.300 ;
        RECT 16.600 106.200 16.900 106.800 ;
        RECT 16.600 105.800 17.000 106.200 ;
        RECT 17.400 103.100 17.800 108.900 ;
        RECT 19.800 108.800 21.000 109.100 ;
        RECT 20.600 105.100 21.000 107.900 ;
        RECT 21.400 105.200 21.700 111.800 ;
        RECT 29.400 109.800 29.800 110.200 ;
        RECT 29.400 109.200 29.700 109.800 ;
        RECT 21.400 104.800 21.800 105.200 ;
        RECT 22.200 103.100 22.600 108.900 ;
        RECT 23.000 106.800 23.400 107.200 ;
        RECT 23.000 106.200 23.300 106.800 ;
        RECT 23.000 105.800 23.400 106.200 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 9.400 96.200 9.700 101.800 ;
        RECT 9.400 95.800 9.800 96.200 ;
        RECT 12.600 95.900 13.000 96.300 ;
        RECT 2.200 94.800 2.600 95.200 ;
        RECT 5.400 95.100 5.800 95.200 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 5.400 94.800 6.600 95.100 ;
        RECT 2.200 94.200 2.500 94.800 ;
        RECT 8.600 94.300 9.000 94.400 ;
        RECT 9.400 94.300 9.800 94.400 ;
        RECT 2.200 93.800 2.600 94.200 ;
        RECT 3.000 93.800 3.400 94.200 ;
        RECT 8.600 94.000 9.800 94.300 ;
        RECT 12.600 94.200 12.900 95.900 ;
        RECT 13.400 95.800 13.800 96.200 ;
        RECT 15.900 95.900 16.300 96.300 ;
        RECT 13.400 95.200 13.700 95.800 ;
        RECT 13.400 94.800 13.800 95.200 ;
        RECT 14.600 94.200 15.000 94.300 ;
        RECT 11.800 93.800 12.200 94.200 ;
        RECT 12.600 93.900 15.000 94.200 ;
        RECT 3.000 93.200 3.300 93.800 ;
        RECT 3.000 92.800 3.400 93.200 ;
        RECT 7.000 92.800 7.400 93.200 ;
        RECT 3.800 86.800 4.200 87.200 ;
        RECT 3.800 85.200 4.100 86.800 ;
        RECT 2.200 84.800 2.600 85.200 ;
        RECT 3.000 85.100 3.400 85.200 ;
        RECT 3.800 85.100 4.200 85.200 ;
        RECT 3.000 84.800 4.200 85.100 ;
        RECT 2.200 84.200 2.500 84.800 ;
        RECT 2.200 83.800 2.600 84.200 ;
        RECT 3.000 83.800 3.400 84.200 ;
        RECT 3.000 83.200 3.300 83.800 ;
        RECT 7.000 83.200 7.300 92.800 ;
        RECT 7.800 91.800 8.200 92.200 ;
        RECT 11.000 91.800 11.400 92.200 ;
        RECT 7.800 86.200 8.100 91.800 ;
        RECT 11.000 89.200 11.300 91.800 ;
        RECT 10.200 88.800 10.600 89.200 ;
        RECT 11.000 88.800 11.400 89.200 ;
        RECT 10.200 88.200 10.500 88.800 ;
        RECT 11.800 88.200 12.100 93.800 ;
        RECT 12.600 93.500 12.900 93.900 ;
        RECT 13.300 93.500 13.700 93.600 ;
        RECT 15.000 93.500 15.400 93.600 ;
        RECT 16.000 93.500 16.300 95.900 ;
        RECT 12.600 93.100 13.000 93.500 ;
        RECT 13.300 93.200 15.400 93.500 ;
        RECT 15.900 93.100 16.300 93.500 ;
        RECT 16.600 93.800 17.000 94.200 ;
        RECT 16.600 89.200 16.900 93.800 ;
        RECT 17.400 93.100 17.800 95.900 ;
        RECT 19.000 92.100 19.400 97.900 ;
        RECT 19.800 95.800 20.200 96.200 ;
        RECT 19.800 95.100 20.100 95.800 ;
        RECT 23.000 95.200 23.300 105.800 ;
        RECT 19.800 94.700 20.200 95.100 ;
        RECT 23.000 94.800 23.400 95.200 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 16.600 88.800 17.000 89.200 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 11.800 87.800 12.200 88.200 ;
        RECT 13.400 88.100 13.800 88.200 ;
        RECT 14.200 88.100 14.600 88.200 ;
        RECT 13.400 87.800 14.600 88.100 ;
        RECT 15.000 88.100 15.400 88.200 ;
        RECT 15.800 88.100 16.200 88.200 ;
        RECT 15.000 87.800 16.200 88.100 ;
        RECT 18.200 88.100 18.600 88.200 ;
        RECT 19.000 88.100 19.400 88.200 ;
        RECT 18.200 87.800 19.400 88.100 ;
        RECT 15.800 86.800 16.200 87.200 ;
        RECT 17.400 86.800 17.800 87.200 ;
        RECT 7.800 85.800 8.200 86.200 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 11.800 86.100 12.200 86.200 ;
        RECT 12.600 86.100 13.000 86.200 ;
        RECT 11.800 85.800 13.000 86.100 ;
        RECT 7.800 84.800 8.200 85.200 ;
        RECT 7.800 84.200 8.100 84.800 ;
        RECT 8.600 84.200 8.900 85.800 ;
        RECT 10.200 85.100 10.600 85.200 ;
        RECT 11.000 85.100 11.400 85.200 ;
        RECT 10.200 84.800 11.400 85.100 ;
        RECT 7.800 83.800 8.200 84.200 ;
        RECT 8.600 83.800 9.000 84.200 ;
        RECT 15.800 83.200 16.100 86.800 ;
        RECT 17.400 85.200 17.700 86.800 ;
        RECT 18.200 86.100 18.600 86.200 ;
        RECT 19.000 86.100 19.400 86.200 ;
        RECT 18.200 85.800 19.400 86.100 ;
        RECT 17.400 84.800 17.800 85.200 ;
        RECT 3.000 82.800 3.400 83.200 ;
        RECT 7.000 82.800 7.400 83.200 ;
        RECT 15.800 82.800 16.200 83.200 ;
        RECT 12.600 81.800 13.000 82.200 ;
        RECT 6.900 75.900 7.300 76.300 ;
        RECT 10.200 75.900 10.600 76.300 ;
        RECT 3.800 74.800 4.200 75.200 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 5.400 75.100 5.800 75.200 ;
        RECT 4.600 74.800 5.800 75.100 ;
        RECT 3.800 74.200 4.100 74.800 ;
        RECT 3.800 73.800 4.200 74.200 ;
        RECT 6.900 73.500 7.200 75.900 ;
        RECT 8.200 74.200 8.600 74.300 ;
        RECT 10.300 74.200 10.600 75.900 ;
        RECT 8.200 73.900 10.600 74.200 ;
        RECT 10.300 73.500 10.600 73.900 ;
        RECT 3.800 72.800 4.200 73.200 ;
        RECT 6.900 73.100 7.300 73.500 ;
        RECT 10.200 73.100 10.600 73.500 ;
        RECT 12.600 73.200 12.900 81.800 ;
        RECT 17.400 76.200 17.700 84.800 ;
        RECT 19.800 81.800 20.200 82.200 ;
        RECT 19.800 77.100 20.100 81.800 ;
        RECT 19.000 76.800 20.100 77.100 ;
        RECT 15.000 75.800 15.400 76.200 ;
        RECT 15.800 75.800 16.200 76.200 ;
        RECT 17.400 75.800 17.800 76.200 ;
        RECT 18.200 75.800 18.600 76.200 ;
        RECT 15.000 75.200 15.300 75.800 ;
        RECT 15.000 74.800 15.400 75.200 ;
        RECT 12.600 72.800 13.000 73.200 ;
        RECT 3.800 72.200 4.100 72.800 ;
        RECT 1.400 72.100 1.800 72.200 ;
        RECT 2.200 72.100 2.600 72.200 ;
        RECT 1.400 71.800 2.600 72.100 ;
        RECT 3.800 71.800 4.200 72.200 ;
        RECT 4.600 71.800 5.000 72.200 ;
        RECT 9.400 71.800 9.800 72.200 ;
        RECT 4.600 69.200 4.900 71.800 ;
        RECT 4.600 68.800 5.000 69.200 ;
        RECT 9.400 68.200 9.700 71.800 ;
        RECT 15.800 69.200 16.100 75.800 ;
        RECT 18.200 74.200 18.500 75.800 ;
        RECT 19.000 75.200 19.300 76.800 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 16.600 73.800 17.000 74.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 16.600 73.200 16.900 73.800 ;
        RECT 16.600 72.800 17.000 73.200 ;
        RECT 19.800 73.100 20.200 75.900 ;
        RECT 20.600 74.200 20.900 93.800 ;
        RECT 23.800 92.100 24.200 97.900 ;
        RECT 24.600 89.200 24.900 105.800 ;
        RECT 27.000 103.100 27.400 108.900 ;
        RECT 29.400 108.800 29.800 109.200 ;
        RECT 30.200 107.200 30.500 124.800 ;
        RECT 33.400 123.100 33.800 128.900 ;
        RECT 34.200 126.800 34.600 127.200 ;
        RECT 35.000 126.800 35.400 127.200 ;
        RECT 37.400 126.800 37.800 127.200 ;
        RECT 34.200 126.300 34.500 126.800 ;
        RECT 34.200 125.900 34.600 126.300 ;
        RECT 31.000 112.100 31.400 117.900 ;
        RECT 31.800 115.800 32.200 116.200 ;
        RECT 31.800 115.100 32.100 115.800 ;
        RECT 35.000 115.200 35.300 126.800 ;
        RECT 37.400 126.200 37.700 126.800 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 38.200 123.100 38.600 128.900 ;
        RECT 43.000 127.800 43.400 128.200 ;
        RECT 53.400 127.800 53.800 128.200 ;
        RECT 43.000 126.200 43.300 127.800 ;
        RECT 51.000 126.800 51.400 127.200 ;
        RECT 41.400 125.800 41.800 126.200 ;
        RECT 43.000 125.800 43.400 126.200 ;
        RECT 47.800 125.800 48.200 126.200 ;
        RECT 41.400 125.200 41.700 125.800 ;
        RECT 47.800 125.200 48.100 125.800 ;
        RECT 41.400 124.800 41.800 125.200 ;
        RECT 43.800 124.800 44.200 125.200 ;
        RECT 47.800 124.800 48.200 125.200 ;
        RECT 43.800 124.200 44.100 124.800 ;
        RECT 43.800 123.800 44.200 124.200 ;
        RECT 46.200 123.800 46.600 124.200 ;
        RECT 45.400 122.800 45.800 123.200 ;
        RECT 39.800 122.100 40.200 122.200 ;
        RECT 40.600 122.100 41.000 122.200 ;
        RECT 39.800 121.800 41.000 122.100 ;
        RECT 42.200 121.800 42.600 122.200 ;
        RECT 31.800 114.700 32.200 115.100 ;
        RECT 35.000 114.800 35.400 115.200 ;
        RECT 35.800 112.100 36.200 117.900 ;
        RECT 39.000 115.100 39.400 115.200 ;
        RECT 39.800 115.100 40.200 115.200 ;
        RECT 39.000 114.800 40.200 115.100 ;
        RECT 39.000 113.100 39.400 113.200 ;
        RECT 39.800 113.100 40.200 113.200 ;
        RECT 39.000 112.800 40.200 113.100 ;
        RECT 40.600 112.800 41.000 113.200 ;
        RECT 40.600 112.200 40.900 112.800 ;
        RECT 38.200 112.100 38.600 112.200 ;
        RECT 39.000 112.100 39.400 112.200 ;
        RECT 38.200 111.800 39.400 112.100 ;
        RECT 40.600 111.800 41.000 112.200 ;
        RECT 42.200 110.200 42.500 121.800 ;
        RECT 45.400 119.200 45.700 122.800 ;
        RECT 45.400 118.800 45.800 119.200 ;
        RECT 43.000 114.800 43.400 115.200 ;
        RECT 44.600 114.800 45.000 115.200 ;
        RECT 43.000 114.200 43.300 114.800 ;
        RECT 44.600 114.200 44.900 114.800 ;
        RECT 43.000 113.800 43.400 114.200 ;
        RECT 44.600 113.800 45.000 114.200 ;
        RECT 43.000 112.800 43.400 113.200 ;
        RECT 43.800 113.100 44.200 113.200 ;
        RECT 44.600 113.100 45.000 113.200 ;
        RECT 43.800 112.800 45.000 113.100 ;
        RECT 43.000 112.200 43.300 112.800 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 42.200 109.800 42.600 110.200 ;
        RECT 35.800 108.800 36.200 109.200 ;
        RECT 40.600 109.100 41.000 109.200 ;
        RECT 41.400 109.100 41.800 109.200 ;
        RECT 40.600 108.800 41.800 109.100 ;
        RECT 43.800 108.800 44.200 109.200 ;
        RECT 31.100 107.800 31.500 107.900 ;
        RECT 31.100 107.500 33.900 107.800 ;
        RECT 34.200 107.500 34.600 107.900 ;
        RECT 30.200 106.800 30.600 107.200 ;
        RECT 31.100 105.100 31.400 107.500 ;
        RECT 31.800 107.400 32.200 107.500 ;
        RECT 33.500 107.400 33.900 107.500 ;
        RECT 34.300 107.100 34.600 107.500 ;
        RECT 31.800 106.800 34.600 107.100 ;
        RECT 35.000 107.800 35.400 108.200 ;
        RECT 35.000 107.200 35.300 107.800 ;
        RECT 35.800 107.200 36.100 108.800 ;
        RECT 43.800 108.200 44.100 108.800 ;
        RECT 39.000 107.500 39.400 107.900 ;
        RECT 42.100 107.800 42.500 107.900 ;
        RECT 43.800 107.800 44.200 108.200 ;
        RECT 39.700 107.500 42.500 107.800 ;
        RECT 35.000 106.800 35.400 107.200 ;
        RECT 35.800 107.100 36.200 107.200 ;
        RECT 36.600 107.100 37.000 107.200 ;
        RECT 35.800 106.800 37.000 107.100 ;
        RECT 37.400 106.800 37.800 107.200 ;
        RECT 39.000 107.100 39.300 107.500 ;
        RECT 39.700 107.400 40.100 107.500 ;
        RECT 41.400 107.400 41.800 107.500 ;
        RECT 39.000 106.800 41.800 107.100 ;
        RECT 31.800 106.100 32.100 106.800 ;
        RECT 31.700 105.700 32.100 106.100 ;
        RECT 34.300 105.100 34.600 106.800 ;
        RECT 37.400 105.200 37.700 106.800 ;
        RECT 31.100 104.700 31.500 105.100 ;
        RECT 34.200 104.700 34.600 105.100 ;
        RECT 35.800 105.100 36.200 105.200 ;
        RECT 36.600 105.100 37.000 105.200 ;
        RECT 35.800 104.800 37.000 105.100 ;
        RECT 37.400 104.800 37.800 105.200 ;
        RECT 39.000 105.100 39.300 106.800 ;
        RECT 41.500 106.100 41.800 106.800 ;
        RECT 41.500 105.700 41.900 106.100 ;
        RECT 42.200 105.100 42.500 107.500 ;
        RECT 46.200 107.200 46.500 123.800 ;
        RECT 51.000 123.200 51.300 126.800 ;
        RECT 52.600 124.800 53.000 125.200 ;
        RECT 52.600 124.200 52.900 124.800 ;
        RECT 52.600 123.800 53.000 124.200 ;
        RECT 53.400 123.200 53.700 127.800 ;
        RECT 55.800 127.500 56.200 127.900 ;
        RECT 56.500 127.500 58.600 127.800 ;
        RECT 59.100 127.500 59.500 127.900 ;
        RECT 55.800 127.100 56.100 127.500 ;
        RECT 56.500 127.400 56.900 127.500 ;
        RECT 58.200 127.400 58.600 127.500 ;
        RECT 55.800 126.800 58.200 127.100 ;
        RECT 55.800 125.100 56.100 126.800 ;
        RECT 57.800 126.700 58.200 126.800 ;
        RECT 58.200 125.800 58.600 126.200 ;
        RECT 55.800 124.700 56.200 125.100 ;
        RECT 58.200 124.200 58.500 125.800 ;
        RECT 59.200 125.100 59.500 127.500 ;
        RECT 59.100 124.700 59.500 125.100 ;
        RECT 59.800 126.800 60.200 127.200 ;
        RECT 59.800 124.200 60.100 126.800 ;
        RECT 60.600 125.100 61.000 127.900 ;
        RECT 61.400 127.800 61.800 128.200 ;
        RECT 61.400 127.200 61.700 127.800 ;
        RECT 61.400 126.800 61.800 127.200 ;
        RECT 58.200 123.800 58.600 124.200 ;
        RECT 59.800 123.800 60.200 124.200 ;
        RECT 51.000 122.800 51.400 123.200 ;
        RECT 53.400 122.800 53.800 123.200 ;
        RECT 62.200 123.100 62.600 128.900 ;
        RECT 63.000 125.900 63.400 126.300 ;
        RECT 63.000 125.200 63.300 125.900 ;
        RECT 66.200 125.800 66.600 126.200 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 51.800 121.800 52.200 122.200 ;
        RECT 51.800 116.200 52.100 121.800 ;
        RECT 51.800 115.800 52.200 116.200 ;
        RECT 52.600 116.100 53.000 116.200 ;
        RECT 53.400 116.100 53.800 116.200 ;
        RECT 52.600 115.800 53.800 116.100 ;
        RECT 54.200 115.800 54.600 116.200 ;
        RECT 55.000 116.100 55.400 116.200 ;
        RECT 55.800 116.100 56.200 116.200 ;
        RECT 55.000 115.800 56.200 116.100 ;
        RECT 58.200 115.800 58.600 116.200 ;
        RECT 54.200 115.200 54.500 115.800 ;
        RECT 58.200 115.200 58.500 115.800 ;
        RECT 47.800 115.100 48.200 115.200 ;
        RECT 48.600 115.100 49.000 115.200 ;
        RECT 47.800 114.800 49.000 115.100 ;
        RECT 54.200 114.800 54.600 115.200 ;
        RECT 58.200 114.800 58.600 115.200 ;
        RECT 59.000 115.100 59.400 115.200 ;
        RECT 59.800 115.100 60.200 115.200 ;
        RECT 59.000 114.800 60.200 115.100 ;
        RECT 47.000 113.800 47.400 114.200 ;
        RECT 50.200 114.100 50.600 114.200 ;
        RECT 51.000 114.100 51.400 114.200 ;
        RECT 50.200 113.800 51.400 114.100 ;
        RECT 54.200 114.100 54.600 114.200 ;
        RECT 55.000 114.100 55.400 114.200 ;
        RECT 54.200 113.800 55.400 114.100 ;
        RECT 55.800 113.800 56.200 114.200 ;
        RECT 56.600 113.800 57.000 114.200 ;
        RECT 47.000 113.200 47.300 113.800 ;
        RECT 55.800 113.200 56.100 113.800 ;
        RECT 56.600 113.200 56.900 113.800 ;
        RECT 47.000 112.800 47.400 113.200 ;
        RECT 55.800 112.800 56.200 113.200 ;
        RECT 56.600 112.800 57.000 113.200 ;
        RECT 60.600 112.800 61.000 113.200 ;
        RECT 61.400 113.100 61.800 113.200 ;
        RECT 62.200 113.100 62.600 113.200 ;
        RECT 63.000 113.100 63.400 115.900 ;
        RECT 61.400 112.800 62.600 113.100 ;
        RECT 50.200 108.800 50.600 109.200 ;
        RECT 50.200 107.200 50.500 108.800 ;
        RECT 51.000 107.500 51.400 107.900 ;
        RECT 51.700 107.500 53.800 107.800 ;
        RECT 54.300 107.500 54.700 107.900 ;
        RECT 43.000 106.800 43.400 107.200 ;
        RECT 46.200 106.800 46.600 107.200 ;
        RECT 47.800 107.100 48.200 107.200 ;
        RECT 48.600 107.100 49.000 107.200 ;
        RECT 47.800 106.800 49.000 107.100 ;
        RECT 50.200 106.800 50.600 107.200 ;
        RECT 51.000 107.100 51.300 107.500 ;
        RECT 51.700 107.400 52.100 107.500 ;
        RECT 53.400 107.400 53.800 107.500 ;
        RECT 51.000 106.800 53.400 107.100 ;
        RECT 43.000 106.200 43.300 106.800 ;
        RECT 43.000 105.800 43.400 106.200 ;
        RECT 44.600 106.100 45.000 106.200 ;
        RECT 45.400 106.100 45.800 106.200 ;
        RECT 44.600 105.800 45.800 106.100 ;
        RECT 46.200 106.100 46.600 106.200 ;
        RECT 47.000 106.100 47.400 106.200 ;
        RECT 46.200 105.800 47.400 106.100 ;
        RECT 27.800 103.800 28.200 104.200 ;
        RECT 26.200 96.800 26.600 97.200 ;
        RECT 26.200 95.200 26.500 96.800 ;
        RECT 26.200 94.800 26.600 95.200 ;
        RECT 27.000 93.100 27.400 95.900 ;
        RECT 27.800 94.200 28.100 103.800 ;
        RECT 32.600 101.800 33.000 102.200 ;
        RECT 27.800 93.800 28.200 94.200 ;
        RECT 28.600 92.100 29.000 97.900 ;
        RECT 30.200 94.800 30.600 95.200 ;
        RECT 30.200 94.200 30.500 94.800 ;
        RECT 30.200 93.800 30.600 94.200 ;
        RECT 31.000 93.800 31.400 94.200 ;
        RECT 21.400 88.800 21.800 89.200 ;
        RECT 24.600 88.800 25.000 89.200 ;
        RECT 21.400 87.200 21.700 88.800 ;
        RECT 23.800 87.500 24.200 87.900 ;
        RECT 24.500 87.500 26.600 87.800 ;
        RECT 27.100 87.500 27.500 87.900 ;
        RECT 21.400 86.800 21.800 87.200 ;
        RECT 23.800 87.100 24.100 87.500 ;
        RECT 24.500 87.400 24.900 87.500 ;
        RECT 26.200 87.400 26.600 87.500 ;
        RECT 23.800 86.800 26.200 87.100 ;
        RECT 21.400 86.200 21.700 86.800 ;
        RECT 21.400 85.800 21.800 86.200 ;
        RECT 23.800 85.100 24.100 86.800 ;
        RECT 25.800 86.700 26.200 86.800 ;
        RECT 27.200 85.100 27.500 87.500 ;
        RECT 23.800 84.700 24.200 85.100 ;
        RECT 27.100 84.700 27.500 85.100 ;
        RECT 27.800 86.800 28.200 87.200 ;
        RECT 27.800 85.200 28.100 86.800 ;
        RECT 27.800 84.800 28.200 85.200 ;
        RECT 28.600 85.100 29.000 87.900 ;
        RECT 27.000 83.800 27.400 84.200 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 20.600 73.200 20.900 73.800 ;
        RECT 20.600 72.800 21.000 73.200 ;
        RECT 17.400 71.800 17.800 72.200 ;
        RECT 21.400 72.100 21.800 77.900 ;
        RECT 26.200 72.100 26.600 77.900 ;
        RECT 17.400 70.200 17.700 71.800 ;
        RECT 21.400 70.800 21.800 71.200 ;
        RECT 17.400 69.800 17.800 70.200 ;
        RECT 21.400 69.200 21.700 70.800 ;
        RECT 27.000 69.200 27.300 83.800 ;
        RECT 30.200 83.100 30.600 88.900 ;
        RECT 31.000 88.200 31.300 93.800 ;
        RECT 31.000 87.800 31.400 88.200 ;
        RECT 31.000 85.900 31.400 86.300 ;
        RECT 31.000 84.200 31.300 85.900 ;
        RECT 31.000 83.800 31.400 84.200 ;
        RECT 28.600 76.800 29.000 77.200 ;
        RECT 28.600 76.200 28.900 76.800 ;
        RECT 28.600 75.800 29.000 76.200 ;
        RECT 29.400 73.100 29.800 75.900 ;
        RECT 31.000 72.100 31.400 77.900 ;
        RECT 32.600 69.200 32.900 101.800 ;
        RECT 37.400 100.200 37.700 104.800 ;
        RECT 39.000 104.700 39.400 105.100 ;
        RECT 42.100 104.700 42.500 105.100 ;
        RECT 44.600 105.100 45.000 105.200 ;
        RECT 45.400 105.100 45.800 105.200 ;
        RECT 44.600 104.800 45.800 105.100 ;
        RECT 51.000 105.100 51.300 106.800 ;
        RECT 53.000 106.700 53.400 106.800 ;
        RECT 53.400 105.800 53.800 106.200 ;
        RECT 51.000 104.700 51.400 105.100 ;
        RECT 53.400 104.200 53.700 105.800 ;
        RECT 54.400 105.100 54.700 107.500 ;
        RECT 54.300 104.700 54.700 105.100 ;
        RECT 55.000 106.800 55.400 107.200 ;
        RECT 53.400 103.800 53.800 104.200 ;
        RECT 54.200 103.800 54.600 104.200 ;
        RECT 35.800 99.800 36.200 100.200 ;
        RECT 37.400 99.800 37.800 100.200 ;
        RECT 35.800 99.200 36.100 99.800 ;
        RECT 54.200 99.200 54.500 103.800 ;
        RECT 35.800 98.800 36.200 99.200 ;
        RECT 54.200 98.800 54.600 99.200 ;
        RECT 55.000 98.100 55.300 106.800 ;
        RECT 55.800 105.100 56.200 107.900 ;
        RECT 56.600 104.200 56.900 112.800 ;
        RECT 56.600 103.800 57.000 104.200 ;
        RECT 57.400 103.100 57.800 108.900 ;
        RECT 58.200 105.900 58.600 106.300 ;
        RECT 58.200 105.200 58.500 105.900 ;
        RECT 58.200 104.800 58.600 105.200 ;
        RECT 33.400 92.100 33.800 97.900 ;
        RECT 40.600 95.800 41.000 96.200 ;
        RECT 40.600 95.200 40.900 95.800 ;
        RECT 38.200 95.100 38.600 95.200 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 38.200 94.800 39.400 95.100 ;
        RECT 40.600 94.800 41.000 95.200 ;
        RECT 38.200 93.800 38.600 94.200 ;
        RECT 40.600 93.800 41.000 94.200 ;
        RECT 38.200 93.200 38.500 93.800 ;
        RECT 40.600 93.200 40.900 93.800 ;
        RECT 36.600 93.100 37.000 93.200 ;
        RECT 37.400 93.100 37.800 93.200 ;
        RECT 36.600 92.800 37.800 93.100 ;
        RECT 38.200 92.800 38.600 93.200 ;
        RECT 40.600 92.800 41.000 93.200 ;
        RECT 41.400 93.100 41.800 95.900 ;
        RECT 36.600 92.100 37.000 92.200 ;
        RECT 37.400 92.100 37.800 92.200 ;
        RECT 36.600 91.800 37.800 92.100 ;
        RECT 37.400 89.100 37.800 89.200 ;
        RECT 38.200 89.100 38.500 92.800 ;
        RECT 43.000 92.100 43.400 97.900 ;
        RECT 43.800 95.800 44.200 96.200 ;
        RECT 43.800 95.100 44.100 95.800 ;
        RECT 46.200 95.100 46.600 95.200 ;
        RECT 47.000 95.100 47.400 95.200 ;
        RECT 43.800 94.700 44.200 95.100 ;
        RECT 46.200 94.800 47.400 95.100 ;
        RECT 47.800 92.100 48.200 97.900 ;
        RECT 54.200 97.800 55.300 98.100 ;
        RECT 52.600 92.800 53.000 93.200 ;
        RECT 52.600 92.200 52.900 92.800 ;
        RECT 50.200 91.800 50.600 92.200 ;
        RECT 52.600 91.800 53.000 92.200 ;
        RECT 50.200 91.200 50.500 91.800 ;
        RECT 50.200 90.800 50.600 91.200 ;
        RECT 35.000 83.100 35.400 88.900 ;
        RECT 37.400 88.800 38.500 89.100 ;
        RECT 38.200 85.100 38.600 87.900 ;
        RECT 39.800 83.100 40.200 88.900 ;
        RECT 43.000 86.800 43.400 87.200 ;
        RECT 43.000 86.200 43.300 86.800 ;
        RECT 43.000 85.800 43.400 86.200 ;
        RECT 36.600 78.800 37.000 79.200 ;
        RECT 34.200 75.100 34.600 75.200 ;
        RECT 35.000 75.100 35.400 75.200 ;
        RECT 34.200 74.800 35.400 75.100 ;
        RECT 35.800 72.100 36.200 77.900 ;
        RECT 35.800 70.800 36.200 71.200 ;
        RECT 12.600 68.800 13.000 69.200 ;
        RECT 15.800 68.800 16.200 69.200 ;
        RECT 21.400 68.800 21.800 69.200 ;
        RECT 27.000 68.800 27.400 69.200 ;
        RECT 32.600 68.800 33.000 69.200 ;
        RECT 12.600 68.200 12.900 68.800 ;
        RECT 2.200 67.800 2.600 68.200 ;
        RECT 2.200 67.200 2.500 67.800 ;
        RECT 3.800 67.500 4.200 67.900 ;
        RECT 7.100 67.500 7.500 67.900 ;
        RECT 2.200 66.800 2.600 67.200 ;
        RECT 3.800 67.100 4.100 67.500 ;
        RECT 3.800 66.800 6.200 67.100 ;
        RECT 3.800 65.100 4.100 66.800 ;
        RECT 5.800 66.700 6.200 66.800 ;
        RECT 7.200 65.100 7.500 67.500 ;
        RECT 8.600 67.800 9.000 68.200 ;
        RECT 9.400 67.800 9.800 68.200 ;
        RECT 12.600 68.100 13.000 68.200 ;
        RECT 12.600 67.800 13.700 68.100 ;
        RECT 8.600 67.200 8.900 67.800 ;
        RECT 8.600 66.800 9.000 67.200 ;
        RECT 10.200 67.100 10.600 67.200 ;
        RECT 11.000 67.100 11.400 67.200 ;
        RECT 10.200 66.800 11.400 67.100 ;
        RECT 13.400 66.200 13.700 67.800 ;
        RECT 15.000 67.800 15.400 68.200 ;
        RECT 17.400 67.800 17.800 68.200 ;
        RECT 15.000 66.200 15.300 67.800 ;
        RECT 17.400 67.200 17.700 67.800 ;
        RECT 19.000 67.500 19.400 67.900 ;
        RECT 22.100 67.800 22.500 67.900 ;
        RECT 19.700 67.500 22.500 67.800 ;
        RECT 15.800 66.800 16.200 67.200 ;
        RECT 17.400 66.800 17.800 67.200 ;
        RECT 19.000 67.100 19.300 67.500 ;
        RECT 19.700 67.400 20.100 67.500 ;
        RECT 21.400 67.400 21.800 67.500 ;
        RECT 19.000 66.800 21.800 67.100 ;
        RECT 15.800 66.200 16.100 66.800 ;
        RECT 13.400 65.800 13.800 66.200 ;
        RECT 15.000 65.800 15.400 66.200 ;
        RECT 15.800 65.800 16.200 66.200 ;
        RECT 3.800 64.700 4.200 65.100 ;
        RECT 7.100 64.700 7.500 65.100 ;
        RECT 15.000 65.100 15.400 65.200 ;
        RECT 15.800 65.100 16.200 65.200 ;
        RECT 15.000 64.800 16.200 65.100 ;
        RECT 19.000 65.100 19.300 66.800 ;
        RECT 21.500 66.100 21.800 66.800 ;
        RECT 21.500 65.700 21.900 66.100 ;
        RECT 22.200 65.100 22.500 67.500 ;
        RECT 24.600 67.500 25.000 67.900 ;
        RECT 27.700 67.800 28.100 67.900 ;
        RECT 25.300 67.500 28.100 67.800 ;
        RECT 19.000 64.700 19.400 65.100 ;
        RECT 22.100 64.700 22.500 65.100 ;
        RECT 23.000 66.800 23.400 67.200 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 24.600 67.100 24.900 67.500 ;
        RECT 25.300 67.400 25.700 67.500 ;
        RECT 27.000 67.400 27.400 67.500 ;
        RECT 24.600 66.800 27.400 67.100 ;
        RECT 23.000 65.200 23.300 66.800 ;
        RECT 23.800 66.200 24.100 66.800 ;
        RECT 23.800 65.800 24.200 66.200 ;
        RECT 23.000 64.800 23.400 65.200 ;
        RECT 24.600 65.100 24.900 66.800 ;
        RECT 27.100 66.100 27.400 66.800 ;
        RECT 27.100 65.700 27.500 66.100 ;
        RECT 27.800 65.100 28.100 67.500 ;
        RECT 28.600 67.800 29.000 68.200 ;
        RECT 28.600 67.200 28.900 67.800 ;
        RECT 30.200 67.500 30.600 67.900 ;
        RECT 33.300 67.800 33.700 67.900 ;
        RECT 30.900 67.500 33.700 67.800 ;
        RECT 28.600 66.800 29.000 67.200 ;
        RECT 29.400 66.800 29.800 67.200 ;
        RECT 30.200 67.100 30.500 67.500 ;
        RECT 30.900 67.400 31.300 67.500 ;
        RECT 32.600 67.400 33.000 67.500 ;
        RECT 30.200 66.800 33.000 67.100 ;
        RECT 24.600 64.700 25.000 65.100 ;
        RECT 27.700 64.700 28.100 65.100 ;
        RECT 29.400 64.200 29.700 66.800 ;
        RECT 30.200 65.100 30.500 66.800 ;
        RECT 31.000 66.100 31.400 66.200 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 31.000 65.800 32.200 66.100 ;
        RECT 32.700 66.100 33.000 66.800 ;
        RECT 32.700 65.700 33.100 66.100 ;
        RECT 33.400 65.100 33.700 67.500 ;
        RECT 30.200 64.700 30.600 65.100 ;
        RECT 33.300 64.700 33.700 65.100 ;
        RECT 35.000 67.800 35.400 68.200 ;
        RECT 19.000 63.800 19.400 64.200 ;
        RECT 29.400 63.800 29.800 64.200 ;
        RECT 5.400 61.800 5.800 62.200 ;
        RECT 12.600 61.800 13.000 62.200 ;
        RECT 1.300 55.900 1.700 56.300 ;
        RECT 1.300 53.500 1.600 55.900 ;
        RECT 3.800 55.800 4.200 56.200 ;
        RECT 4.600 55.900 5.000 56.300 ;
        RECT 3.800 55.200 4.100 55.800 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 2.600 54.200 3.000 54.300 ;
        RECT 4.700 54.200 5.000 55.900 ;
        RECT 2.600 53.900 5.000 54.200 ;
        RECT 2.200 53.500 2.600 53.600 ;
        RECT 3.900 53.500 4.300 53.600 ;
        RECT 4.700 53.500 5.000 53.900 ;
        RECT 5.400 54.200 5.700 61.800 ;
        RECT 12.600 59.200 12.900 61.800 ;
        RECT 19.000 59.200 19.300 63.800 ;
        RECT 11.000 58.800 11.400 59.200 ;
        RECT 12.600 58.800 13.000 59.200 ;
        RECT 19.000 58.800 19.400 59.200 ;
        RECT 31.000 59.100 31.400 59.200 ;
        RECT 31.800 59.100 32.200 59.200 ;
        RECT 31.000 58.800 32.200 59.100 ;
        RECT 5.400 53.800 5.800 54.200 ;
        RECT 1.300 53.100 1.700 53.500 ;
        RECT 2.200 53.200 4.300 53.500 ;
        RECT 3.000 52.800 3.400 53.200 ;
        RECT 4.600 53.100 5.000 53.500 ;
        RECT 6.200 53.100 6.600 55.900 ;
        RECT 7.800 52.100 8.200 57.900 ;
        RECT 8.600 55.800 9.000 56.200 ;
        RECT 8.600 55.100 8.900 55.800 ;
        RECT 8.600 54.700 9.000 55.100 ;
        RECT 8.600 52.800 9.000 53.200 ;
        RECT 8.600 49.200 8.900 52.800 ;
        RECT 8.600 48.800 9.000 49.200 ;
        RECT 3.800 47.500 4.200 47.900 ;
        RECT 7.100 47.500 7.500 47.900 ;
        RECT 3.800 47.100 4.100 47.500 ;
        RECT 3.800 46.800 6.200 47.100 ;
        RECT 3.000 45.800 3.400 46.200 ;
        RECT 3.000 45.200 3.300 45.800 ;
        RECT 3.000 44.800 3.400 45.200 ;
        RECT 3.800 45.100 4.100 46.800 ;
        RECT 5.800 46.700 6.200 46.800 ;
        RECT 6.200 45.800 6.600 46.200 ;
        RECT 3.800 44.700 4.200 45.100 ;
        RECT 6.200 44.200 6.500 45.800 ;
        RECT 7.200 45.100 7.500 47.500 ;
        RECT 11.000 47.200 11.300 58.800 ;
        RECT 11.800 54.800 12.200 55.200 ;
        RECT 11.800 52.200 12.100 54.800 ;
        RECT 11.800 51.800 12.200 52.200 ;
        RECT 12.600 52.100 13.000 57.900 ;
        RECT 24.600 56.800 25.000 57.200 ;
        RECT 16.500 55.900 16.900 56.300 ;
        RECT 19.800 55.900 20.200 56.300 ;
        RECT 24.600 56.200 24.900 56.800 ;
        RECT 35.000 56.200 35.300 67.800 ;
        RECT 16.500 53.500 16.800 55.900 ;
        RECT 17.800 54.200 18.200 54.300 ;
        RECT 19.900 54.200 20.200 55.900 ;
        RECT 23.800 55.800 24.200 56.200 ;
        RECT 24.600 55.800 25.000 56.200 ;
        RECT 29.400 55.800 29.800 56.200 ;
        RECT 35.000 55.800 35.400 56.200 ;
        RECT 23.800 55.200 24.100 55.800 ;
        RECT 29.400 55.200 29.700 55.800 ;
        RECT 23.800 54.800 24.200 55.200 ;
        RECT 26.200 55.100 26.600 55.200 ;
        RECT 27.000 55.100 27.400 55.200 ;
        RECT 26.200 54.800 27.400 55.100 ;
        RECT 29.400 54.800 29.800 55.200 ;
        RECT 32.600 54.800 33.000 55.200 ;
        RECT 32.600 54.200 32.900 54.800 ;
        RECT 17.800 53.900 20.200 54.200 ;
        RECT 17.400 53.500 17.800 53.600 ;
        RECT 19.100 53.500 19.500 53.600 ;
        RECT 19.900 53.500 20.200 53.900 ;
        RECT 15.000 52.800 15.400 53.200 ;
        RECT 16.500 53.100 16.900 53.500 ;
        RECT 17.400 53.200 19.500 53.500 ;
        RECT 17.400 52.800 17.800 53.200 ;
        RECT 19.800 53.100 20.200 53.500 ;
        RECT 20.600 53.800 21.000 54.200 ;
        RECT 21.400 53.800 21.800 54.200 ;
        RECT 32.600 53.800 33.000 54.200 ;
        RECT 15.000 52.200 15.300 52.800 ;
        RECT 15.000 51.800 15.400 52.200 ;
        RECT 18.200 51.800 18.600 52.200 ;
        RECT 12.600 47.500 13.000 47.900 ;
        RECT 15.700 47.800 16.100 47.900 ;
        RECT 13.300 47.500 16.100 47.800 ;
        RECT 11.000 46.800 11.400 47.200 ;
        RECT 12.600 47.100 12.900 47.500 ;
        RECT 13.300 47.400 13.700 47.500 ;
        RECT 15.000 47.400 15.400 47.500 ;
        RECT 12.600 46.800 15.400 47.100 ;
        RECT 9.400 46.100 9.800 46.200 ;
        RECT 10.200 46.100 10.600 46.200 ;
        RECT 9.400 45.800 10.600 46.100 ;
        RECT 7.100 44.700 7.500 45.100 ;
        RECT 7.800 45.100 8.200 45.200 ;
        RECT 8.600 45.100 9.000 45.200 ;
        RECT 7.800 44.800 9.000 45.100 ;
        RECT 12.600 45.100 12.900 46.800 ;
        RECT 13.400 46.100 13.800 46.200 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 13.400 45.800 14.600 46.100 ;
        RECT 15.100 46.100 15.400 46.800 ;
        RECT 15.100 45.700 15.500 46.100 ;
        RECT 15.800 45.100 16.100 47.500 ;
        RECT 16.600 47.800 17.000 48.200 ;
        RECT 16.600 47.200 16.900 47.800 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 17.400 45.100 17.800 47.900 ;
        RECT 18.200 47.200 18.500 51.800 ;
        RECT 18.200 46.800 18.600 47.200 ;
        RECT 12.600 44.700 13.000 45.100 ;
        RECT 15.700 44.700 16.100 45.100 ;
        RECT 6.200 43.800 6.600 44.200 ;
        RECT 19.000 43.100 19.400 48.900 ;
        RECT 19.800 45.900 20.200 46.300 ;
        RECT 19.800 45.200 20.100 45.900 ;
        RECT 19.800 44.800 20.200 45.200 ;
        RECT 18.200 41.800 18.600 42.200 ;
        RECT 7.000 36.800 7.400 37.200 ;
        RECT 1.500 35.900 1.900 36.300 ;
        RECT 4.600 35.900 5.000 36.300 ;
        RECT 1.500 33.500 1.800 35.900 ;
        RECT 2.100 34.900 2.500 35.300 ;
        RECT 2.200 34.200 2.500 34.900 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 3.000 34.800 4.200 35.100 ;
        RECT 4.700 34.200 5.000 35.900 ;
        RECT 7.000 36.200 7.300 36.800 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 9.400 36.100 9.800 36.200 ;
        RECT 10.200 36.100 10.600 36.200 ;
        RECT 9.400 35.800 10.600 36.100 ;
        RECT 14.200 35.900 14.600 36.300 ;
        RECT 15.800 36.100 16.200 36.200 ;
        RECT 16.600 36.100 17.000 36.200 ;
        RECT 11.000 35.100 11.400 35.200 ;
        RECT 11.800 35.100 12.200 35.200 ;
        RECT 11.000 34.800 12.200 35.100 ;
        RECT 12.600 34.800 13.000 35.200 ;
        RECT 2.200 33.900 5.000 34.200 ;
        RECT 2.200 33.500 2.600 33.600 ;
        RECT 3.900 33.500 4.300 33.600 ;
        RECT 4.700 33.500 5.000 33.900 ;
        RECT 12.600 34.200 12.900 34.800 ;
        RECT 14.200 34.200 14.500 35.900 ;
        RECT 15.800 35.800 17.000 36.100 ;
        RECT 17.300 35.900 17.700 36.300 ;
        RECT 16.700 34.900 17.100 35.300 ;
        RECT 16.700 34.200 17.000 34.900 ;
        RECT 12.600 33.800 13.000 34.200 ;
        RECT 14.200 33.900 17.000 34.200 ;
        RECT 1.500 33.200 4.300 33.500 ;
        RECT 1.500 33.100 1.900 33.200 ;
        RECT 4.600 33.100 5.000 33.500 ;
        RECT 14.200 33.500 14.500 33.900 ;
        RECT 14.900 33.500 15.300 33.600 ;
        RECT 16.600 33.500 17.000 33.600 ;
        RECT 17.400 33.500 17.700 35.900 ;
        RECT 18.200 35.200 18.500 41.800 ;
        RECT 20.600 39.200 20.900 53.800 ;
        RECT 21.400 53.200 21.700 53.800 ;
        RECT 21.400 52.800 21.800 53.200 ;
        RECT 24.600 53.100 25.000 53.200 ;
        RECT 25.400 53.100 25.800 53.200 ;
        RECT 24.600 52.800 25.800 53.100 ;
        RECT 26.200 52.800 26.600 53.200 ;
        RECT 26.200 49.200 26.500 52.800 ;
        RECT 23.000 46.800 23.400 47.200 ;
        RECT 23.000 46.200 23.300 46.800 ;
        RECT 23.000 45.800 23.400 46.200 ;
        RECT 23.800 43.100 24.200 48.900 ;
        RECT 26.200 48.800 26.600 49.200 ;
        RECT 35.800 48.200 36.100 70.800 ;
        RECT 36.600 66.200 36.900 78.800 ;
        RECT 37.400 74.100 37.800 74.200 ;
        RECT 38.200 74.100 38.600 74.200 ;
        RECT 37.400 73.800 38.600 74.100 ;
        RECT 39.000 73.100 39.400 75.900 ;
        RECT 40.600 72.100 41.000 77.900 ;
        RECT 41.400 75.800 41.800 76.200 ;
        RECT 41.400 75.100 41.700 75.800 ;
        RECT 43.000 75.200 43.300 85.800 ;
        RECT 44.600 83.100 45.000 88.900 ;
        RECT 47.800 86.100 48.200 86.200 ;
        RECT 48.600 86.100 49.000 86.200 ;
        RECT 47.800 85.800 49.000 86.100 ;
        RECT 49.400 85.100 49.800 87.900 ;
        RECT 50.200 87.800 50.600 88.200 ;
        RECT 50.200 87.200 50.500 87.800 ;
        RECT 50.200 86.800 50.600 87.200 ;
        RECT 51.000 83.100 51.400 88.900 ;
        RECT 51.800 85.900 52.200 86.300 ;
        RECT 51.800 85.200 52.100 85.900 ;
        RECT 51.800 84.800 52.200 85.200 ;
        RECT 41.400 74.700 41.800 75.100 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 43.000 74.200 43.300 74.800 ;
        RECT 43.000 73.800 43.400 74.200 ;
        RECT 36.600 65.800 37.000 66.200 ;
        RECT 37.400 65.100 37.800 67.900 ;
        RECT 39.000 63.100 39.400 68.900 ;
        RECT 39.800 68.800 40.200 69.200 ;
        RECT 39.800 66.300 40.100 68.800 ;
        RECT 43.000 67.200 43.300 73.800 ;
        RECT 45.400 72.100 45.800 77.900 ;
        RECT 50.200 73.100 50.600 75.900 ;
        RECT 47.800 72.100 48.200 72.200 ;
        RECT 48.600 72.100 49.000 72.200 ;
        RECT 51.800 72.100 52.200 77.900 ;
        RECT 52.600 74.700 53.000 75.100 ;
        RECT 52.600 74.200 52.900 74.700 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 52.600 72.800 53.000 73.200 ;
        RECT 47.800 71.800 49.000 72.100 ;
        RECT 43.000 66.800 43.400 67.200 ;
        RECT 39.800 65.900 40.200 66.300 ;
        RECT 43.000 66.200 43.300 66.800 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 39.000 53.100 39.400 55.900 ;
        RECT 39.800 54.800 40.200 55.200 ;
        RECT 39.800 54.200 40.100 54.800 ;
        RECT 39.800 53.800 40.200 54.200 ;
        RECT 40.600 52.100 41.000 57.900 ;
        RECT 42.200 54.800 42.600 55.200 ;
        RECT 42.200 54.200 42.500 54.800 ;
        RECT 43.000 54.200 43.300 65.800 ;
        RECT 43.800 63.100 44.200 68.900 ;
        RECT 48.600 65.100 49.000 67.900 ;
        RECT 49.400 67.800 49.800 68.200 ;
        RECT 49.400 67.200 49.700 67.800 ;
        RECT 49.400 66.800 49.800 67.200 ;
        RECT 47.800 62.800 48.200 63.200 ;
        RECT 50.200 63.100 50.600 68.900 ;
        RECT 52.600 67.200 52.900 72.800 ;
        RECT 52.600 66.800 53.000 67.200 ;
        RECT 51.000 65.900 51.400 66.300 ;
        RECT 51.000 65.200 51.300 65.900 ;
        RECT 51.000 64.800 51.400 65.200 ;
        RECT 46.200 61.800 46.600 62.200 ;
        RECT 42.200 53.800 42.600 54.200 ;
        RECT 43.000 53.800 43.400 54.200 ;
        RECT 43.800 51.800 44.200 52.200 ;
        RECT 45.400 52.100 45.800 57.900 ;
        RECT 46.200 52.200 46.500 61.800 ;
        RECT 47.800 59.200 48.100 62.800 ;
        RECT 52.600 60.800 53.000 61.200 ;
        RECT 52.600 59.200 52.900 60.800 ;
        RECT 47.800 58.800 48.200 59.200 ;
        RECT 52.600 58.800 53.000 59.200 ;
        RECT 54.200 58.200 54.500 97.800 ;
        RECT 60.600 97.200 60.900 112.800 ;
        RECT 64.600 112.100 65.000 117.900 ;
        RECT 65.400 115.800 65.800 116.200 ;
        RECT 65.400 115.100 65.700 115.800 ;
        RECT 65.400 114.700 65.800 115.100 ;
        RECT 66.200 114.200 66.500 125.800 ;
        RECT 67.000 123.100 67.400 128.900 ;
        RECT 107.000 128.800 107.400 129.200 ;
        RECT 107.000 128.200 107.300 128.800 ;
        RECT 71.000 127.500 71.400 127.900 ;
        RECT 71.700 127.500 73.800 127.800 ;
        RECT 74.300 127.500 74.700 127.900 ;
        RECT 70.200 126.800 70.600 127.200 ;
        RECT 71.000 127.100 71.300 127.500 ;
        RECT 71.700 127.400 72.100 127.500 ;
        RECT 73.400 127.400 73.800 127.500 ;
        RECT 71.000 126.800 73.400 127.100 ;
        RECT 69.400 121.800 69.800 122.200 ;
        RECT 69.400 121.200 69.700 121.800 ;
        RECT 69.400 120.800 69.800 121.200 ;
        RECT 67.800 114.800 68.200 115.200 ;
        RECT 66.200 113.800 66.600 114.200 ;
        RECT 61.400 105.800 61.800 106.200 ;
        RECT 61.400 105.200 61.700 105.800 ;
        RECT 61.400 104.800 61.800 105.200 ;
        RECT 62.200 103.100 62.600 108.900 ;
        RECT 65.400 105.100 65.800 107.900 ;
        RECT 66.200 107.200 66.500 113.800 ;
        RECT 66.200 106.800 66.600 107.200 ;
        RECT 66.200 106.200 66.500 106.800 ;
        RECT 66.200 105.800 66.600 106.200 ;
        RECT 66.200 103.800 66.600 104.200 ;
        RECT 64.600 102.100 65.000 102.200 ;
        RECT 65.400 102.100 65.800 102.200 ;
        RECT 64.600 101.800 65.800 102.100 ;
        RECT 60.600 96.800 61.000 97.200 ;
        RECT 60.600 96.200 60.900 96.800 ;
        RECT 58.200 95.800 58.600 96.200 ;
        RECT 59.800 95.800 60.200 96.200 ;
        RECT 60.600 95.800 61.000 96.200 ;
        RECT 58.200 94.200 58.500 95.800 ;
        RECT 59.000 94.800 59.400 95.200 ;
        RECT 56.600 93.800 57.000 94.200 ;
        RECT 58.200 93.800 58.600 94.200 ;
        RECT 56.600 93.200 56.900 93.800 ;
        RECT 59.000 93.200 59.300 94.800 ;
        RECT 55.000 93.100 55.400 93.200 ;
        RECT 55.800 93.100 56.200 93.200 ;
        RECT 55.000 92.800 56.200 93.100 ;
        RECT 56.600 92.800 57.000 93.200 ;
        RECT 59.000 93.100 59.400 93.200 ;
        RECT 59.800 93.100 60.100 95.800 ;
        RECT 66.200 95.200 66.500 103.800 ;
        RECT 67.000 103.100 67.400 108.900 ;
        RECT 67.000 101.800 67.400 102.200 ;
        RECT 60.600 94.800 61.000 95.200 ;
        RECT 66.200 94.800 66.600 95.200 ;
        RECT 60.600 94.200 60.900 94.800 ;
        RECT 60.600 93.800 61.000 94.200 ;
        RECT 63.000 94.100 63.400 94.200 ;
        RECT 63.800 94.100 64.200 94.200 ;
        RECT 63.000 93.800 64.200 94.100 ;
        RECT 64.600 93.800 65.000 94.200 ;
        RECT 64.600 93.200 64.900 93.800 ;
        RECT 59.000 92.800 60.100 93.100 ;
        RECT 63.000 93.100 63.400 93.200 ;
        RECT 63.800 93.100 64.200 93.200 ;
        RECT 63.000 92.800 64.200 93.100 ;
        RECT 64.600 92.800 65.000 93.200 ;
        RECT 55.800 83.100 56.200 88.900 ;
        RECT 56.600 82.100 56.900 92.800 ;
        RECT 55.800 81.800 56.900 82.100 ;
        RECT 57.400 91.800 57.800 92.200 ;
        RECT 61.400 91.800 61.800 92.200 ;
        RECT 63.000 91.800 63.400 92.200 ;
        RECT 57.400 88.200 57.700 91.800 ;
        RECT 57.400 87.800 57.800 88.200 ;
        RECT 58.200 88.100 58.600 88.200 ;
        RECT 59.000 88.100 59.400 88.200 ;
        RECT 58.200 87.800 59.400 88.100 ;
        RECT 55.000 63.100 55.400 68.900 ;
        RECT 55.000 61.800 55.400 62.200 ;
        RECT 55.000 59.200 55.300 61.800 ;
        RECT 55.800 59.200 56.100 81.800 ;
        RECT 57.400 79.200 57.700 87.800 ;
        RECT 61.400 86.200 61.700 91.800 ;
        RECT 63.000 89.200 63.300 91.800 ;
        RECT 63.000 88.800 63.400 89.200 ;
        RECT 63.800 86.800 64.200 87.200 ;
        RECT 61.400 85.800 61.800 86.200 ;
        RECT 63.800 82.200 64.100 86.800 ;
        RECT 58.200 82.100 58.600 82.200 ;
        RECT 59.000 82.100 59.400 82.200 ;
        RECT 58.200 81.800 59.400 82.100 ;
        RECT 63.800 81.800 64.200 82.200 ;
        RECT 57.400 78.800 57.800 79.200 ;
        RECT 56.600 72.100 57.000 77.900 ;
        RECT 57.400 77.800 57.800 78.200 ;
        RECT 63.800 77.800 64.200 78.200 ;
        RECT 57.400 69.200 57.700 77.800 ;
        RECT 63.800 77.200 64.100 77.800 ;
        RECT 64.600 77.200 64.900 92.800 ;
        RECT 66.200 90.200 66.500 94.800 ;
        RECT 66.200 89.800 66.600 90.200 ;
        RECT 67.000 89.200 67.300 101.800 ;
        RECT 67.800 99.200 68.100 114.800 ;
        RECT 69.400 112.100 69.800 117.900 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 68.600 105.200 68.900 105.800 ;
        RECT 68.600 104.800 69.000 105.200 ;
        RECT 70.200 102.200 70.500 126.800 ;
        RECT 71.000 125.100 71.300 126.800 ;
        RECT 73.000 126.700 73.400 126.800 ;
        RECT 74.400 125.100 74.700 127.500 ;
        RECT 76.500 127.500 76.900 127.900 ;
        RECT 77.400 127.500 79.500 127.800 ;
        RECT 79.800 127.500 80.200 127.900 ;
        RECT 71.000 124.700 71.400 125.100 ;
        RECT 74.300 124.700 74.700 125.100 ;
        RECT 75.800 126.800 76.200 127.200 ;
        RECT 75.800 124.200 76.100 126.800 ;
        RECT 76.500 125.100 76.800 127.500 ;
        RECT 77.400 127.400 77.800 127.500 ;
        RECT 79.100 127.400 79.500 127.500 ;
        RECT 79.900 127.100 80.200 127.500 ;
        RECT 83.800 127.500 84.200 127.900 ;
        RECT 84.500 127.500 86.600 127.800 ;
        RECT 87.100 127.500 87.500 127.900 ;
        RECT 77.800 126.800 80.200 127.100 ;
        RECT 80.600 127.100 81.000 127.200 ;
        RECT 81.400 127.100 81.800 127.200 ;
        RECT 80.600 126.800 81.800 127.100 ;
        RECT 83.800 127.100 84.100 127.500 ;
        RECT 84.500 127.400 84.900 127.500 ;
        RECT 86.200 127.400 86.600 127.500 ;
        RECT 83.800 126.800 86.200 127.100 ;
        RECT 77.800 126.700 78.200 126.800 ;
        RECT 79.000 125.800 79.400 126.200 ;
        RECT 79.000 125.200 79.300 125.800 ;
        RECT 76.500 124.700 76.900 125.100 ;
        RECT 79.000 124.800 79.400 125.200 ;
        RECT 79.900 125.100 80.200 126.800 ;
        RECT 79.800 124.700 80.200 125.100 ;
        RECT 83.800 125.100 84.100 126.800 ;
        RECT 85.800 126.700 86.200 126.800 ;
        RECT 86.200 125.800 86.600 126.200 ;
        RECT 83.800 124.700 84.200 125.100 ;
        RECT 86.200 124.200 86.500 125.800 ;
        RECT 87.200 125.100 87.500 127.500 ;
        RECT 106.200 127.800 106.600 128.200 ;
        RECT 107.000 127.800 107.400 128.200 ;
        RECT 109.400 127.800 109.800 128.200 ;
        RECT 106.200 127.200 106.500 127.800 ;
        RECT 109.400 127.200 109.700 127.800 ;
        RECT 113.400 127.500 113.800 127.900 ;
        RECT 114.100 127.500 116.200 127.800 ;
        RECT 116.700 127.500 117.100 127.900 ;
        RECT 87.100 124.700 87.500 125.100 ;
        RECT 87.800 126.800 88.200 127.200 ;
        RECT 93.400 126.800 93.800 127.200 ;
        RECT 94.200 126.800 94.600 127.200 ;
        RECT 98.200 126.800 98.600 127.200 ;
        RECT 100.600 126.800 101.000 127.200 ;
        RECT 106.200 126.800 106.600 127.200 ;
        RECT 107.800 126.800 108.200 127.200 ;
        RECT 109.400 126.800 109.800 127.200 ;
        RECT 112.600 126.800 113.000 127.200 ;
        RECT 113.400 127.100 113.700 127.500 ;
        RECT 114.100 127.400 114.500 127.500 ;
        RECT 115.800 127.400 116.200 127.500 ;
        RECT 113.400 126.800 115.800 127.100 ;
        RECT 75.800 123.800 76.200 124.200 ;
        RECT 86.200 123.800 86.600 124.200 ;
        RECT 72.600 123.100 73.000 123.200 ;
        RECT 73.400 123.100 73.800 123.200 ;
        RECT 72.600 122.800 73.800 123.100 ;
        RECT 75.800 119.200 76.100 123.800 ;
        RECT 79.000 121.800 79.400 122.200 ;
        RECT 79.000 119.200 79.300 121.800 ;
        RECT 87.800 120.200 88.100 126.800 ;
        RECT 93.400 126.200 93.700 126.800 ;
        RECT 88.600 125.800 89.000 126.200 ;
        RECT 89.400 125.800 89.800 126.200 ;
        RECT 90.200 125.800 90.600 126.200 ;
        RECT 91.800 126.100 92.200 126.200 ;
        RECT 92.600 126.100 93.000 126.200 ;
        RECT 91.800 125.800 93.000 126.100 ;
        RECT 93.400 125.800 93.800 126.200 ;
        RECT 88.600 125.200 88.900 125.800 ;
        RECT 88.600 124.800 89.000 125.200 ;
        RECT 89.400 123.100 89.700 125.800 ;
        RECT 90.200 124.200 90.500 125.800 ;
        RECT 91.800 124.800 92.200 125.200 ;
        RECT 91.800 124.200 92.100 124.800 ;
        RECT 90.200 123.800 90.600 124.200 ;
        RECT 91.800 123.800 92.200 124.200 ;
        RECT 89.400 122.800 90.500 123.100 ;
        RECT 87.800 119.800 88.200 120.200 ;
        RECT 90.200 119.200 90.500 122.800 ;
        RECT 94.200 122.200 94.500 126.800 ;
        RECT 96.600 126.100 97.000 126.200 ;
        RECT 96.600 125.800 97.700 126.100 ;
        RECT 95.800 123.800 96.200 124.200 ;
        RECT 95.800 123.200 96.100 123.800 ;
        RECT 95.800 122.800 96.200 123.200 ;
        RECT 96.600 122.800 97.000 123.200 ;
        RECT 96.600 122.200 96.900 122.800 ;
        RECT 91.000 121.800 91.400 122.200 ;
        RECT 94.200 121.800 94.600 122.200 ;
        RECT 96.600 121.800 97.000 122.200 ;
        RECT 75.800 118.800 76.200 119.200 ;
        RECT 79.000 118.800 79.400 119.200 ;
        RECT 90.200 118.800 90.600 119.200 ;
        RECT 91.000 117.200 91.300 121.800 ;
        RECT 92.600 119.800 93.000 120.200 ;
        RECT 86.200 116.800 86.600 117.200 ;
        RECT 89.400 117.100 89.800 117.200 ;
        RECT 90.200 117.100 90.600 117.200 ;
        RECT 89.400 116.800 90.600 117.100 ;
        RECT 91.000 116.800 91.400 117.200 ;
        RECT 73.300 115.900 73.700 116.300 ;
        RECT 76.600 115.900 77.000 116.300 ;
        RECT 73.300 113.500 73.600 115.900 ;
        RECT 74.600 114.200 75.000 114.300 ;
        RECT 76.700 114.200 77.000 115.900 ;
        RECT 81.400 115.800 81.800 116.200 ;
        RECT 81.400 114.200 81.700 115.800 ;
        RECT 86.200 115.200 86.500 116.800 ;
        RECT 90.200 116.200 90.500 116.800 ;
        RECT 87.000 116.100 87.400 116.200 ;
        RECT 87.800 116.100 88.200 116.200 ;
        RECT 87.000 115.800 88.900 116.100 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 85.400 114.200 85.700 114.800 ;
        RECT 74.600 113.900 77.000 114.200 ;
        RECT 74.200 113.500 74.600 113.600 ;
        RECT 75.900 113.500 76.300 113.600 ;
        RECT 76.700 113.500 77.000 113.900 ;
        RECT 79.000 114.100 79.400 114.200 ;
        RECT 79.000 113.800 80.100 114.100 ;
        RECT 73.300 113.100 73.700 113.500 ;
        RECT 74.200 113.200 76.300 113.500 ;
        RECT 71.800 112.100 72.200 112.200 ;
        RECT 72.600 112.100 73.000 112.200 ;
        RECT 71.800 111.800 73.000 112.100 ;
        RECT 71.800 103.100 72.200 108.900 ;
        RECT 75.000 107.200 75.300 113.200 ;
        RECT 76.600 113.100 77.000 113.500 ;
        RECT 78.200 110.800 78.600 111.200 ;
        RECT 78.200 109.200 78.500 110.800 ;
        RECT 78.200 108.800 78.600 109.200 ;
        RECT 75.900 107.800 76.300 107.900 ;
        RECT 75.900 107.500 78.700 107.800 ;
        RECT 79.000 107.500 79.400 107.900 ;
        RECT 75.000 106.800 75.400 107.200 ;
        RECT 75.000 104.200 75.300 106.800 ;
        RECT 75.900 105.100 76.200 107.500 ;
        RECT 76.600 107.400 77.000 107.500 ;
        RECT 78.300 107.400 78.700 107.500 ;
        RECT 79.100 107.100 79.400 107.500 ;
        RECT 76.600 106.800 79.400 107.100 ;
        RECT 76.600 106.100 76.900 106.800 ;
        RECT 76.500 105.700 76.900 106.100 ;
        RECT 77.400 105.800 77.800 106.200 ;
        RECT 75.900 104.700 76.300 105.100 ;
        RECT 75.000 103.800 75.400 104.200 ;
        RECT 70.200 101.800 70.600 102.200 ;
        RECT 74.200 101.800 74.600 102.200 ;
        RECT 67.800 98.800 68.200 99.200 ;
        RECT 74.200 98.200 74.500 101.800 ;
        RECT 74.200 97.800 74.600 98.200 ;
        RECT 71.800 95.800 72.200 96.200 ;
        RECT 75.000 96.100 75.400 96.200 ;
        RECT 75.800 96.100 76.200 96.200 ;
        RECT 75.000 95.800 76.200 96.100 ;
        RECT 76.600 95.800 77.000 96.200 ;
        RECT 67.800 94.800 68.200 95.200 ;
        RECT 68.600 94.800 69.000 95.200 ;
        RECT 70.200 95.100 70.600 95.200 ;
        RECT 71.000 95.100 71.400 95.200 ;
        RECT 70.200 94.800 71.400 95.100 ;
        RECT 67.800 93.200 68.100 94.800 ;
        RECT 68.600 94.200 68.900 94.800 ;
        RECT 68.600 93.800 69.000 94.200 ;
        RECT 69.400 94.100 69.800 94.200 ;
        RECT 70.200 94.100 70.600 94.200 ;
        RECT 69.400 93.800 70.600 94.100 ;
        RECT 71.800 93.200 72.100 95.800 ;
        RECT 72.600 94.800 73.000 95.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 75.000 94.800 75.400 95.200 ;
        RECT 72.600 94.200 72.900 94.800 ;
        RECT 72.600 93.800 73.000 94.200 ;
        RECT 67.800 92.800 68.200 93.200 ;
        RECT 71.800 92.800 72.200 93.200 ;
        RECT 67.800 89.200 68.100 92.800 ;
        RECT 71.800 91.800 72.200 92.200 ;
        RECT 71.800 91.200 72.100 91.800 ;
        RECT 71.800 90.800 72.200 91.200 ;
        RECT 73.400 91.100 73.700 94.800 ;
        RECT 75.000 94.200 75.300 94.800 ;
        RECT 75.000 93.800 75.400 94.200 ;
        RECT 76.600 93.200 76.900 95.800 ;
        RECT 75.800 93.100 76.200 93.200 ;
        RECT 76.600 93.100 77.000 93.200 ;
        RECT 75.800 92.800 77.000 93.100 ;
        RECT 77.400 92.100 77.700 105.800 ;
        RECT 79.100 105.100 79.400 106.800 ;
        RECT 79.800 107.200 80.100 113.800 ;
        RECT 81.400 113.800 81.800 114.200 ;
        RECT 84.600 113.800 85.000 114.200 ;
        RECT 85.400 113.800 85.800 114.200 ;
        RECT 81.400 109.200 81.700 113.800 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 81.400 108.800 81.800 109.200 ;
        RECT 79.800 106.800 80.200 107.200 ;
        RECT 80.600 107.100 81.000 107.200 ;
        RECT 81.400 107.100 81.800 107.200 ;
        RECT 80.600 106.800 81.800 107.100 ;
        RECT 79.800 106.200 80.100 106.800 ;
        RECT 79.800 105.800 80.200 106.200 ;
        RECT 79.000 104.700 79.400 105.100 ;
        RECT 82.200 105.200 82.500 111.800 ;
        RECT 84.600 109.200 84.900 113.800 ;
        RECT 88.600 113.200 88.900 115.800 ;
        RECT 89.400 115.800 89.800 116.200 ;
        RECT 90.200 115.800 90.600 116.200 ;
        RECT 88.600 112.800 89.000 113.200 ;
        RECT 87.800 111.800 88.200 112.200 ;
        RECT 84.600 108.800 85.000 109.200 ;
        RECT 87.800 108.200 88.100 111.800 ;
        RECT 89.400 111.200 89.700 115.800 ;
        RECT 90.200 114.800 90.600 115.200 ;
        RECT 90.200 114.200 90.500 114.800 ;
        RECT 90.200 113.800 90.600 114.200 ;
        RECT 89.400 110.800 89.800 111.200 ;
        RECT 90.200 109.200 90.500 113.800 ;
        RECT 92.600 113.200 92.900 119.800 ;
        RECT 94.200 119.200 94.500 121.800 ;
        RECT 97.400 121.200 97.700 125.800 ;
        RECT 98.200 125.200 98.500 126.800 ;
        RECT 98.200 124.800 98.600 125.200 ;
        RECT 95.800 120.800 96.200 121.200 ;
        RECT 97.400 120.800 97.800 121.200 ;
        RECT 95.800 119.200 96.100 120.800 ;
        RECT 98.200 120.200 98.500 124.800 ;
        RECT 98.200 119.800 98.600 120.200 ;
        RECT 100.600 119.200 100.900 126.800 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 104.600 125.800 105.000 126.200 ;
        RECT 107.000 125.800 107.400 126.200 ;
        RECT 93.400 118.800 93.800 119.200 ;
        RECT 94.200 118.800 94.600 119.200 ;
        RECT 95.800 118.800 96.200 119.200 ;
        RECT 100.600 118.800 101.000 119.200 ;
        RECT 93.400 118.200 93.700 118.800 ;
        RECT 93.400 117.800 93.800 118.200 ;
        RECT 95.000 117.800 95.400 118.200 ;
        RECT 95.000 117.200 95.300 117.800 ;
        RECT 95.000 116.800 95.400 117.200 ;
        RECT 95.800 115.800 96.200 116.200 ;
        RECT 96.600 115.800 97.000 116.200 ;
        RECT 99.000 115.800 99.400 116.200 ;
        RECT 95.800 115.200 96.100 115.800 ;
        RECT 95.800 114.800 96.200 115.200 ;
        RECT 96.600 114.200 96.900 115.800 ;
        RECT 99.000 114.200 99.300 115.800 ;
        RECT 99.800 114.800 100.200 115.200 ;
        RECT 96.600 113.800 97.000 114.200 ;
        RECT 97.400 114.100 97.800 114.200 ;
        RECT 98.200 114.100 98.600 114.200 ;
        RECT 97.400 113.800 98.600 114.100 ;
        RECT 99.000 113.800 99.400 114.200 ;
        RECT 99.800 113.200 100.100 114.800 ;
        RECT 92.600 112.800 93.000 113.200 ;
        RECT 97.400 112.800 97.800 113.200 ;
        RECT 99.800 112.800 100.200 113.200 ;
        RECT 92.600 109.200 92.900 112.800 ;
        RECT 93.400 111.800 93.800 112.200 ;
        RECT 93.400 109.200 93.700 111.800 ;
        RECT 97.400 111.200 97.700 112.800 ;
        RECT 101.400 112.200 101.700 125.800 ;
        RECT 104.600 119.200 104.900 125.800 ;
        RECT 106.200 123.800 106.600 124.200 ;
        RECT 104.600 118.800 105.000 119.200 ;
        RECT 104.600 117.800 105.000 118.200 ;
        RECT 104.600 113.200 104.900 117.800 ;
        RECT 106.200 113.200 106.500 123.800 ;
        RECT 107.000 119.200 107.300 125.800 ;
        RECT 107.000 118.800 107.400 119.200 ;
        RECT 107.000 115.200 107.300 118.800 ;
        RECT 107.000 114.800 107.400 115.200 ;
        RECT 107.800 114.200 108.100 126.800 ;
        RECT 112.600 126.200 112.900 126.800 ;
        RECT 109.400 126.100 109.800 126.200 ;
        RECT 110.200 126.100 110.600 126.200 ;
        RECT 109.400 125.800 110.600 126.100 ;
        RECT 111.000 125.800 111.400 126.200 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 112.600 125.800 113.000 126.200 ;
        RECT 111.000 121.200 111.300 125.800 ;
        RECT 111.800 125.200 112.100 125.800 ;
        RECT 111.800 124.800 112.200 125.200 ;
        RECT 113.400 125.100 113.700 126.800 ;
        RECT 115.400 126.700 115.800 126.800 ;
        RECT 116.800 125.100 117.100 127.500 ;
        RECT 117.400 127.800 117.800 128.200 ;
        RECT 120.600 127.800 121.000 128.200 ;
        RECT 121.400 127.800 121.800 128.200 ;
        RECT 117.400 127.200 117.700 127.800 ;
        RECT 117.400 126.800 117.800 127.200 ;
        RECT 119.000 126.800 119.400 127.200 ;
        RECT 113.400 124.700 113.800 125.100 ;
        RECT 116.700 124.700 117.100 125.100 ;
        RECT 118.200 125.800 118.600 126.200 ;
        RECT 114.200 121.800 114.600 122.200 ;
        RECT 111.000 120.800 111.400 121.200 ;
        RECT 112.600 118.800 113.000 119.200 ;
        RECT 112.600 118.200 112.900 118.800 ;
        RECT 112.600 117.800 113.000 118.200 ;
        RECT 114.200 116.200 114.500 121.800 ;
        RECT 118.200 117.200 118.500 125.800 ;
        RECT 119.000 118.200 119.300 126.800 ;
        RECT 119.000 117.800 119.400 118.200 ;
        RECT 118.200 116.800 118.600 117.200 ;
        RECT 114.200 115.800 114.600 116.200 ;
        RECT 115.700 115.900 116.100 116.300 ;
        RECT 119.000 115.900 119.400 116.300 ;
        RECT 112.600 114.800 113.000 115.200 ;
        RECT 112.600 114.200 112.900 114.800 ;
        RECT 107.000 113.800 107.400 114.200 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 112.600 113.800 113.000 114.200 ;
        RECT 115.000 113.800 115.400 114.200 ;
        RECT 104.600 112.800 105.000 113.200 ;
        RECT 106.200 112.800 106.600 113.200 ;
        RECT 107.000 112.200 107.300 113.800 ;
        RECT 101.400 111.800 101.800 112.200 ;
        RECT 107.000 111.800 107.400 112.200 ;
        RECT 97.400 110.800 97.800 111.200 ;
        RECT 90.200 108.800 90.600 109.200 ;
        RECT 92.600 108.800 93.000 109.200 ;
        RECT 93.400 108.800 93.800 109.200 ;
        RECT 101.400 108.800 101.800 109.200 ;
        RECT 85.400 107.800 85.800 108.200 ;
        RECT 87.800 107.800 88.200 108.200 ;
        RECT 91.800 108.100 92.200 108.200 ;
        RECT 92.600 108.100 93.000 108.200 ;
        RECT 98.200 108.100 98.600 108.200 ;
        RECT 91.800 107.800 93.000 108.100 ;
        RECT 97.400 107.800 98.600 108.100 ;
        RECT 83.800 106.800 84.200 107.200 ;
        RECT 83.800 106.200 84.100 106.800 ;
        RECT 83.000 105.800 83.400 106.200 ;
        RECT 83.800 105.800 84.200 106.200 ;
        RECT 82.200 104.800 82.600 105.200 ;
        RECT 82.200 102.200 82.500 104.800 ;
        RECT 82.200 101.800 82.600 102.200 ;
        RECT 83.000 101.200 83.300 105.800 ;
        RECT 83.000 100.800 83.400 101.200 ;
        RECT 83.800 98.200 84.100 105.800 ;
        RECT 85.400 104.200 85.700 107.800 ;
        RECT 87.000 106.100 87.400 106.200 ;
        RECT 87.800 106.100 88.200 106.200 ;
        RECT 87.000 105.800 88.200 106.100 ;
        RECT 91.000 105.800 91.400 106.200 ;
        RECT 88.600 105.100 89.000 105.200 ;
        RECT 89.400 105.100 89.800 105.200 ;
        RECT 88.600 104.800 89.800 105.100 ;
        RECT 85.400 103.800 85.800 104.200 ;
        RECT 88.600 104.100 89.000 104.200 ;
        RECT 88.600 103.800 89.700 104.100 ;
        RECT 87.800 103.100 88.200 103.200 ;
        RECT 88.600 103.100 89.000 103.200 ;
        RECT 87.800 102.800 89.000 103.100 ;
        RECT 87.000 99.800 87.400 100.200 ;
        RECT 87.000 99.200 87.300 99.800 ;
        RECT 89.400 99.200 89.700 103.800 ;
        RECT 90.200 103.800 90.600 104.200 ;
        RECT 91.000 104.100 91.300 105.800 ;
        RECT 91.800 105.200 92.100 107.800 ;
        RECT 94.200 106.800 94.600 107.200 ;
        RECT 95.000 106.800 95.400 107.200 ;
        RECT 96.600 106.800 97.000 107.200 ;
        RECT 91.800 104.800 92.200 105.200 ;
        RECT 91.000 103.800 92.100 104.100 ;
        RECT 90.200 103.200 90.500 103.800 ;
        RECT 90.200 102.800 90.600 103.200 ;
        RECT 91.800 99.200 92.100 103.800 ;
        RECT 94.200 103.200 94.500 106.800 ;
        RECT 95.000 106.200 95.300 106.800 ;
        RECT 95.000 105.800 95.400 106.200 ;
        RECT 95.800 105.800 96.200 106.200 ;
        RECT 95.800 105.200 96.100 105.800 ;
        RECT 96.600 105.200 96.900 106.800 ;
        RECT 95.800 104.800 96.200 105.200 ;
        RECT 96.600 104.800 97.000 105.200 ;
        RECT 94.200 102.800 94.600 103.200 ;
        RECT 96.600 102.200 96.900 104.800 ;
        RECT 97.400 104.200 97.700 107.800 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 99.000 106.800 99.400 107.200 ;
        RECT 98.200 106.200 98.500 106.800 ;
        RECT 99.000 106.200 99.300 106.800 ;
        RECT 98.200 105.800 98.600 106.200 ;
        RECT 99.000 105.800 99.400 106.200 ;
        RECT 97.400 103.800 97.800 104.200 ;
        RECT 96.600 101.800 97.000 102.200 ;
        RECT 97.400 99.200 97.700 103.800 ;
        RECT 99.800 101.800 100.200 102.200 ;
        RECT 84.600 99.100 85.000 99.200 ;
        RECT 85.400 99.100 85.800 99.200 ;
        RECT 84.600 98.800 85.800 99.100 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 89.400 98.800 89.800 99.200 ;
        RECT 91.800 98.800 92.200 99.200 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 99.800 98.200 100.100 101.800 ;
        RECT 101.400 99.200 101.700 108.800 ;
        RECT 115.000 108.200 115.300 113.800 ;
        RECT 115.700 113.500 116.000 115.900 ;
        RECT 117.000 114.200 117.400 114.300 ;
        RECT 119.100 114.200 119.400 115.900 ;
        RECT 120.600 116.200 120.900 127.800 ;
        RECT 121.400 127.200 121.700 127.800 ;
        RECT 127.000 127.500 127.400 127.900 ;
        RECT 127.700 127.500 129.800 127.800 ;
        RECT 130.300 127.500 130.700 127.900 ;
        RECT 121.400 126.800 121.800 127.200 ;
        RECT 126.200 126.800 126.600 127.200 ;
        RECT 127.000 127.100 127.300 127.500 ;
        RECT 127.700 127.400 128.100 127.500 ;
        RECT 129.400 127.400 129.800 127.500 ;
        RECT 127.000 126.800 129.400 127.100 ;
        RECT 121.400 126.100 121.800 126.200 ;
        RECT 122.200 126.100 122.600 126.200 ;
        RECT 121.400 125.800 122.600 126.100 ;
        RECT 123.800 125.800 124.200 126.200 ;
        RECT 123.000 124.800 123.400 125.200 ;
        RECT 123.000 119.200 123.300 124.800 ;
        RECT 123.800 123.200 124.100 125.800 ;
        RECT 126.200 125.200 126.500 126.800 ;
        RECT 126.200 124.800 126.600 125.200 ;
        RECT 127.000 125.100 127.300 126.800 ;
        RECT 129.000 126.700 129.400 126.800 ;
        RECT 130.400 125.100 130.700 127.500 ;
        RECT 135.000 127.800 135.400 128.200 ;
        RECT 135.800 127.800 136.200 128.200 ;
        RECT 147.000 128.100 147.400 128.200 ;
        RECT 147.800 128.100 148.200 128.200 ;
        RECT 127.000 124.700 127.400 125.100 ;
        RECT 130.300 124.700 130.700 125.100 ;
        RECT 131.000 126.800 131.400 127.200 ;
        RECT 131.000 124.200 131.300 126.800 ;
        RECT 135.000 126.200 135.300 127.800 ;
        RECT 135.800 127.200 136.100 127.800 ;
        RECT 142.200 127.500 142.600 127.900 ;
        RECT 145.300 127.800 145.700 127.900 ;
        RECT 147.000 127.800 148.200 128.100 ;
        RECT 142.900 127.500 145.700 127.800 ;
        RECT 135.800 126.800 136.200 127.200 ;
        RECT 136.600 126.800 137.000 127.200 ;
        RECT 137.400 127.100 137.800 127.200 ;
        RECT 138.200 127.100 138.600 127.200 ;
        RECT 137.400 126.800 138.600 127.100 ;
        RECT 141.400 126.800 141.800 127.200 ;
        RECT 142.200 127.100 142.500 127.500 ;
        RECT 142.900 127.400 143.300 127.500 ;
        RECT 144.600 127.400 145.000 127.500 ;
        RECT 142.200 126.800 145.000 127.100 ;
        RECT 131.800 125.800 132.200 126.200 ;
        RECT 132.600 125.800 133.000 126.200 ;
        RECT 135.000 125.800 135.400 126.200 ;
        RECT 131.800 125.200 132.100 125.800 ;
        RECT 131.800 124.800 132.200 125.200 ;
        RECT 124.600 124.100 125.000 124.200 ;
        RECT 125.400 124.100 125.800 124.200 ;
        RECT 124.600 123.800 125.800 124.100 ;
        RECT 127.800 124.100 128.200 124.200 ;
        RECT 128.600 124.100 129.000 124.200 ;
        RECT 127.800 123.800 129.000 124.100 ;
        RECT 131.000 123.800 131.400 124.200 ;
        RECT 123.800 122.800 124.200 123.200 ;
        RECT 132.600 122.200 132.900 125.800 ;
        RECT 133.400 123.800 133.800 124.200 ;
        RECT 125.400 121.800 125.800 122.200 ;
        RECT 132.600 121.800 133.000 122.200 ;
        RECT 125.400 119.200 125.700 121.800 ;
        RECT 133.400 121.200 133.700 123.800 ;
        RECT 134.200 123.100 134.600 123.200 ;
        RECT 135.000 123.100 135.400 123.200 ;
        RECT 134.200 122.800 135.400 123.100 ;
        RECT 136.600 121.200 136.900 126.800 ;
        RECT 137.400 125.800 137.800 126.200 ;
        RECT 139.000 125.800 139.400 126.200 ;
        RECT 139.800 125.800 140.200 126.200 ;
        RECT 137.400 122.200 137.700 125.800 ;
        RECT 139.000 125.200 139.300 125.800 ;
        RECT 139.000 124.800 139.400 125.200 ;
        RECT 138.200 123.800 138.600 124.200 ;
        RECT 137.400 121.800 137.800 122.200 ;
        RECT 133.400 120.800 133.800 121.200 ;
        RECT 136.600 120.800 137.000 121.200 ;
        RECT 135.000 119.800 135.400 120.200 ;
        RECT 123.000 118.800 123.400 119.200 ;
        RECT 125.400 118.800 125.800 119.200 ;
        RECT 122.200 117.800 122.600 118.200 ;
        RECT 124.600 117.800 125.000 118.200 ;
        RECT 127.800 117.800 128.200 118.200 ;
        RECT 122.200 117.200 122.500 117.800 ;
        RECT 124.600 117.200 124.900 117.800 ;
        RECT 121.400 116.800 121.800 117.200 ;
        RECT 122.200 116.800 122.600 117.200 ;
        RECT 124.600 116.800 125.000 117.200 ;
        RECT 126.200 116.800 126.600 117.200 ;
        RECT 120.600 115.800 121.000 116.200 ;
        RECT 121.400 115.200 121.700 116.800 ;
        RECT 126.200 116.200 126.500 116.800 ;
        RECT 126.200 115.800 126.600 116.200 ;
        RECT 121.400 114.800 121.800 115.200 ;
        RECT 125.400 114.800 125.800 115.200 ;
        RECT 117.000 113.900 119.400 114.200 ;
        RECT 116.600 113.500 117.000 113.600 ;
        RECT 118.300 113.500 118.700 113.600 ;
        RECT 119.100 113.500 119.400 113.900 ;
        RECT 115.700 113.100 116.100 113.500 ;
        RECT 116.600 113.200 118.700 113.500 ;
        RECT 118.200 112.200 118.500 113.200 ;
        RECT 119.000 113.100 119.400 113.500 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 123.800 114.100 124.200 114.200 ;
        RECT 124.600 114.100 125.000 114.200 ;
        RECT 123.800 113.800 125.000 114.100 ;
        RECT 119.800 113.200 120.100 113.800 ;
        RECT 125.400 113.200 125.700 114.800 ;
        RECT 127.800 114.200 128.100 117.800 ;
        RECT 131.000 115.900 131.400 116.300 ;
        RECT 134.100 115.900 134.500 116.300 ;
        RECT 131.000 114.200 131.300 115.900 ;
        RECT 133.500 114.900 133.900 115.300 ;
        RECT 133.500 114.200 133.800 114.900 ;
        RECT 127.800 113.800 128.200 114.200 ;
        RECT 130.200 113.800 130.600 114.200 ;
        RECT 131.000 113.900 133.800 114.200 ;
        RECT 119.800 112.800 120.200 113.200 ;
        RECT 125.400 112.800 125.800 113.200 ;
        RECT 128.600 113.100 129.000 113.200 ;
        RECT 129.400 113.100 129.800 113.200 ;
        RECT 128.600 112.800 129.800 113.100 ;
        RECT 118.200 111.800 118.600 112.200 ;
        RECT 109.400 107.800 109.800 108.200 ;
        RECT 115.000 107.800 115.400 108.200 ;
        RECT 123.000 107.800 123.400 108.200 ;
        RECT 107.000 106.800 107.400 107.200 ;
        RECT 107.000 106.200 107.300 106.800 ;
        RECT 109.400 106.200 109.700 107.800 ;
        RECT 112.600 107.100 113.000 107.200 ;
        RECT 113.400 107.100 113.800 107.200 ;
        RECT 112.600 106.800 113.800 107.100 ;
        RECT 121.400 106.800 121.800 107.200 ;
        RECT 104.600 105.800 105.000 106.200 ;
        RECT 107.000 105.800 107.400 106.200 ;
        RECT 107.800 105.800 108.200 106.200 ;
        RECT 109.400 105.800 109.800 106.200 ;
        RECT 115.000 106.100 115.400 106.200 ;
        RECT 118.200 106.100 118.600 106.200 ;
        RECT 119.000 106.100 119.400 106.200 ;
        RECT 115.000 105.800 116.100 106.100 ;
        RECT 118.200 105.800 119.400 106.100 ;
        RECT 119.800 106.100 120.200 106.200 ;
        RECT 120.600 106.100 121.000 106.200 ;
        RECT 119.800 105.800 121.000 106.100 ;
        RECT 104.600 105.200 104.900 105.800 ;
        RECT 107.800 105.200 108.100 105.800 ;
        RECT 102.200 104.800 102.600 105.200 ;
        RECT 104.600 104.800 105.000 105.200 ;
        RECT 105.400 104.800 105.800 105.200 ;
        RECT 107.800 104.800 108.200 105.200 ;
        RECT 108.600 104.800 109.000 105.200 ;
        RECT 111.000 104.800 111.400 105.200 ;
        RECT 111.800 104.800 112.200 105.200 ;
        RECT 115.000 104.800 115.400 105.200 ;
        RECT 101.400 98.800 101.800 99.200 ;
        RECT 83.800 97.800 84.200 98.200 ;
        RECT 95.800 97.800 96.200 98.200 ;
        RECT 99.800 97.800 100.200 98.200 ;
        RECT 79.000 97.100 79.400 97.200 ;
        RECT 79.800 97.100 80.200 97.200 ;
        RECT 79.000 96.800 80.200 97.100 ;
        RECT 85.400 96.800 85.800 97.200 ;
        RECT 87.000 96.800 87.400 97.200 ;
        RECT 92.600 97.100 93.000 97.200 ;
        RECT 93.400 97.100 93.800 97.200 ;
        RECT 92.600 96.800 93.800 97.100 ;
        RECT 94.200 96.800 94.600 97.200 ;
        RECT 85.400 96.200 85.700 96.800 ;
        RECT 82.200 96.100 82.600 96.200 ;
        RECT 83.000 96.100 83.400 96.200 ;
        RECT 82.200 95.800 83.400 96.100 ;
        RECT 85.400 95.800 85.800 96.200 ;
        RECT 72.600 90.800 73.700 91.100 ;
        RECT 76.600 91.800 77.700 92.100 ;
        RECT 79.800 94.800 80.200 95.200 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 83.800 95.100 84.200 95.200 ;
        RECT 83.000 94.800 84.200 95.100 ;
        RECT 68.600 89.800 69.000 90.200 ;
        RECT 68.600 89.200 68.900 89.800 ;
        RECT 72.600 89.200 72.900 90.800 ;
        RECT 76.600 89.200 76.900 91.800 ;
        RECT 65.400 88.800 65.800 89.200 ;
        RECT 67.000 88.800 67.400 89.200 ;
        RECT 67.800 88.800 68.200 89.200 ;
        RECT 68.600 88.800 69.000 89.200 ;
        RECT 72.600 88.800 73.000 89.200 ;
        RECT 75.800 88.800 76.200 89.200 ;
        RECT 76.600 88.800 77.000 89.200 ;
        RECT 65.400 88.200 65.700 88.800 ;
        RECT 65.400 87.800 65.800 88.200 ;
        RECT 65.400 87.100 65.800 87.200 ;
        RECT 66.200 87.100 66.600 87.200 ;
        RECT 65.400 86.800 66.600 87.100 ;
        RECT 67.800 86.800 68.200 87.200 ;
        RECT 71.800 86.800 72.200 87.200 ;
        RECT 73.400 86.800 73.800 87.200 ;
        RECT 67.800 85.200 68.100 86.800 ;
        RECT 71.800 86.200 72.100 86.800 ;
        RECT 71.000 85.800 71.400 86.200 ;
        RECT 71.800 85.800 72.200 86.200 ;
        RECT 71.000 85.200 71.300 85.800 ;
        RECT 66.200 84.800 66.600 85.200 ;
        RECT 67.800 84.800 68.200 85.200 ;
        RECT 68.600 84.800 69.000 85.200 ;
        RECT 71.000 84.800 71.400 85.200 ;
        RECT 58.200 77.100 58.600 77.200 ;
        RECT 59.000 77.100 59.400 77.200 ;
        RECT 58.200 76.800 59.400 77.100 ;
        RECT 59.800 77.100 60.200 77.200 ;
        RECT 60.600 77.100 61.000 77.200 ;
        RECT 59.800 76.800 61.000 77.100 ;
        RECT 62.200 77.100 62.600 77.200 ;
        RECT 63.000 77.100 63.400 77.200 ;
        RECT 62.200 76.800 63.400 77.100 ;
        RECT 63.800 76.800 64.200 77.200 ;
        RECT 64.600 76.800 65.000 77.200 ;
        RECT 61.400 76.100 61.800 76.200 ;
        RECT 62.200 76.100 62.600 76.200 ;
        RECT 61.400 75.800 62.600 76.100 ;
        RECT 59.800 74.100 60.200 74.200 ;
        RECT 59.000 73.800 60.200 74.100 ;
        RECT 59.000 72.200 59.300 73.800 ;
        RECT 63.000 73.200 63.300 76.800 ;
        RECT 64.600 75.800 65.000 76.200 ;
        RECT 64.600 75.200 64.900 75.800 ;
        RECT 63.800 74.800 64.200 75.200 ;
        RECT 64.600 74.800 65.000 75.200 ;
        RECT 63.800 74.200 64.100 74.800 ;
        RECT 66.200 74.200 66.500 84.800 ;
        RECT 67.800 76.200 68.100 84.800 ;
        RECT 68.600 84.200 68.900 84.800 ;
        RECT 68.600 83.800 69.000 84.200 ;
        RECT 68.600 77.200 68.900 83.800 ;
        RECT 68.600 76.800 69.000 77.200 ;
        RECT 67.800 75.800 68.200 76.200 ;
        RECT 70.200 75.800 70.600 76.200 ;
        RECT 67.000 75.100 67.400 75.200 ;
        RECT 67.800 75.100 68.200 75.200 ;
        RECT 67.000 74.800 68.200 75.100 ;
        RECT 63.800 73.800 64.200 74.200 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 67.000 74.100 67.400 74.200 ;
        RECT 66.200 73.800 67.400 74.100 ;
        RECT 63.000 72.800 63.400 73.200 ;
        RECT 59.000 71.800 59.400 72.200 ;
        RECT 59.800 71.800 60.200 72.200 ;
        RECT 63.800 72.100 64.100 73.800 ;
        RECT 64.600 73.100 65.000 73.200 ;
        RECT 65.400 73.100 65.800 73.200 ;
        RECT 64.600 72.800 65.800 73.100 ;
        RECT 63.000 71.800 64.100 72.100 ;
        RECT 66.200 71.800 66.600 72.200 ;
        RECT 59.000 71.200 59.300 71.800 ;
        RECT 59.000 70.800 59.400 71.200 ;
        RECT 57.400 68.800 57.800 69.200 ;
        RECT 58.200 66.800 58.600 67.200 ;
        RECT 58.200 60.200 58.500 66.800 ;
        RECT 58.200 59.800 58.600 60.200 ;
        RECT 55.000 58.800 55.400 59.200 ;
        RECT 55.800 58.800 56.200 59.200 ;
        RECT 47.800 57.800 48.200 58.200 ;
        RECT 54.200 57.800 54.600 58.200 ;
        RECT 46.200 51.800 46.600 52.200 ;
        RECT 43.000 48.800 43.400 49.200 ;
        RECT 43.000 48.200 43.300 48.800 ;
        RECT 43.800 48.200 44.100 51.800 ;
        RECT 47.800 49.200 48.100 57.800 ;
        RECT 59.000 57.200 59.300 70.800 ;
        RECT 59.800 69.200 60.100 71.800 ;
        RECT 59.800 68.800 60.200 69.200 ;
        RECT 60.600 68.800 61.000 69.200 ;
        RECT 60.600 67.200 60.900 68.800 ;
        RECT 60.600 66.800 61.000 67.200 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 62.200 66.200 62.500 66.800 ;
        RECT 62.200 65.800 62.600 66.200 ;
        RECT 60.600 64.800 61.000 65.200 ;
        RECT 61.400 65.100 61.800 65.200 ;
        RECT 62.200 65.100 62.600 65.200 ;
        RECT 61.400 64.800 62.600 65.100 ;
        RECT 50.200 56.800 50.600 57.200 ;
        RECT 55.800 56.800 56.200 57.200 ;
        RECT 59.000 56.800 59.400 57.200 ;
        RECT 50.200 55.200 50.500 56.800 ;
        RECT 55.800 56.200 56.100 56.800 ;
        RECT 60.600 56.200 60.900 64.800 ;
        RECT 63.000 57.200 63.300 71.800 ;
        RECT 66.200 68.200 66.500 71.800 ;
        RECT 66.200 67.800 66.600 68.200 ;
        RECT 67.800 68.100 68.200 68.200 ;
        RECT 67.800 67.800 68.900 68.100 ;
        RECT 68.600 67.200 68.900 67.800 ;
        RECT 69.400 67.800 69.800 68.200 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 67.800 66.800 68.200 67.200 ;
        RECT 68.600 66.800 69.000 67.200 ;
        RECT 64.600 66.200 64.900 66.800 ;
        RECT 67.800 66.200 68.100 66.800 ;
        RECT 69.400 66.200 69.700 67.800 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 67.800 65.800 68.200 66.200 ;
        RECT 69.400 65.800 69.800 66.200 ;
        RECT 65.400 65.200 65.700 65.800 ;
        RECT 64.600 64.800 65.000 65.200 ;
        RECT 65.400 64.800 65.800 65.200 ;
        RECT 63.800 63.800 64.200 64.200 ;
        RECT 63.800 62.200 64.100 63.800 ;
        RECT 64.600 63.200 64.900 64.800 ;
        RECT 67.000 63.800 67.400 64.200 ;
        RECT 64.600 62.800 65.000 63.200 ;
        RECT 67.000 62.200 67.300 63.800 ;
        RECT 70.200 63.200 70.500 75.800 ;
        RECT 71.000 75.200 71.300 84.800 ;
        RECT 73.400 84.200 73.700 86.800 ;
        RECT 74.200 85.800 74.600 86.200 ;
        RECT 73.400 83.800 73.800 84.200 ;
        RECT 74.200 83.100 74.500 85.800 ;
        RECT 73.400 82.800 74.500 83.100 ;
        RECT 72.600 76.800 73.000 77.200 ;
        RECT 71.800 75.800 72.200 76.200 ;
        RECT 71.800 75.200 72.100 75.800 ;
        RECT 71.000 74.800 71.400 75.200 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 72.600 74.200 72.900 76.800 ;
        RECT 73.400 75.200 73.700 82.800 ;
        RECT 75.800 79.200 76.100 88.800 ;
        RECT 77.400 86.800 77.800 87.200 ;
        RECT 77.400 86.200 77.700 86.800 ;
        RECT 77.400 85.800 77.800 86.200 ;
        RECT 76.600 84.800 77.000 85.200 ;
        RECT 79.000 84.800 79.400 85.200 ;
        RECT 76.600 84.200 76.900 84.800 ;
        RECT 76.600 83.800 77.000 84.200 ;
        RECT 75.800 78.800 76.200 79.200 ;
        RECT 79.000 77.200 79.300 84.800 ;
        RECT 79.000 76.800 79.400 77.200 ;
        RECT 79.800 76.200 80.100 94.800 ;
        RECT 80.600 93.800 81.000 94.200 ;
        RECT 83.000 94.100 83.400 94.200 ;
        RECT 83.800 94.100 84.200 94.200 ;
        RECT 83.000 93.800 84.200 94.100 ;
        RECT 86.200 93.800 86.600 94.200 ;
        RECT 80.600 89.200 80.900 93.800 ;
        RECT 84.600 91.800 85.000 92.200 ;
        RECT 80.600 88.800 81.000 89.200 ;
        RECT 83.800 87.800 84.200 88.200 ;
        RECT 83.800 87.200 84.100 87.800 ;
        RECT 80.600 87.100 81.000 87.200 ;
        RECT 81.400 87.100 81.800 87.200 ;
        RECT 80.600 86.800 81.800 87.100 ;
        RECT 82.200 87.100 82.600 87.200 ;
        RECT 83.000 87.100 83.400 87.200 ;
        RECT 82.200 86.800 83.400 87.100 ;
        RECT 83.800 86.800 84.200 87.200 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 82.200 85.200 82.500 85.800 ;
        RECT 82.200 84.800 82.600 85.200 ;
        RECT 83.800 76.200 84.100 86.800 ;
        RECT 84.600 86.200 84.900 91.800 ;
        RECT 86.200 91.200 86.500 93.800 ;
        RECT 86.200 90.800 86.600 91.200 ;
        RECT 86.200 89.800 86.600 90.200 ;
        RECT 86.200 89.200 86.500 89.800 ;
        RECT 86.200 88.800 86.600 89.200 ;
        RECT 87.000 88.200 87.300 96.800 ;
        RECT 94.200 96.200 94.500 96.800 ;
        RECT 95.800 96.200 96.100 97.800 ;
        RECT 101.400 96.800 101.800 97.200 ;
        RECT 87.800 95.800 88.200 96.200 ;
        RECT 88.600 96.100 89.000 96.200 ;
        RECT 89.400 96.100 89.800 96.200 ;
        RECT 88.600 95.800 89.800 96.100 ;
        RECT 94.200 95.800 94.600 96.200 ;
        RECT 95.800 96.100 96.200 96.200 ;
        RECT 96.600 96.100 97.000 96.200 ;
        RECT 95.800 95.800 97.000 96.100 ;
        RECT 98.200 96.100 98.600 96.200 ;
        RECT 99.000 96.100 99.400 96.200 ;
        RECT 98.200 95.800 99.400 96.100 ;
        RECT 87.800 95.200 88.100 95.800 ;
        RECT 101.400 95.200 101.700 96.800 ;
        RECT 87.800 94.800 88.200 95.200 ;
        RECT 91.800 94.800 92.200 95.200 ;
        RECT 93.400 94.800 93.800 95.200 ;
        RECT 101.400 94.800 101.800 95.200 ;
        RECT 90.200 93.800 90.600 94.200 ;
        RECT 90.200 92.200 90.500 93.800 ;
        RECT 91.800 92.200 92.100 94.800 ;
        RECT 90.200 91.800 90.600 92.200 ;
        RECT 91.800 91.800 92.200 92.200 ;
        RECT 90.200 90.800 90.600 91.200 ;
        RECT 90.200 88.200 90.500 90.800 ;
        RECT 91.800 89.200 92.100 91.800 ;
        RECT 91.800 88.800 92.200 89.200 ;
        RECT 86.200 87.800 86.600 88.200 ;
        RECT 87.000 87.800 87.400 88.200 ;
        RECT 90.200 87.800 90.600 88.200 ;
        RECT 84.600 85.800 85.000 86.200 ;
        RECT 84.600 78.200 84.900 85.800 ;
        RECT 84.600 77.800 85.000 78.200 ;
        RECT 85.400 76.800 85.800 77.200 ;
        RECT 85.400 76.200 85.700 76.800 ;
        RECT 79.800 75.800 80.200 76.200 ;
        RECT 83.800 75.800 84.200 76.200 ;
        RECT 85.400 75.800 85.800 76.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 74.200 75.100 74.600 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 74.200 74.800 75.400 75.100 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 77.400 75.100 77.800 75.200 ;
        RECT 76.600 74.800 77.800 75.100 ;
        RECT 79.800 75.100 80.200 75.200 ;
        RECT 80.600 75.100 81.000 75.200 ;
        RECT 79.800 74.800 81.000 75.100 ;
        RECT 72.600 73.800 73.000 74.200 ;
        RECT 71.000 72.800 71.400 73.200 ;
        RECT 70.200 62.800 70.600 63.200 ;
        RECT 63.800 61.800 64.200 62.200 ;
        RECT 67.000 61.800 67.400 62.200 ;
        RECT 70.200 59.800 70.600 60.200 ;
        RECT 70.200 59.200 70.500 59.800 ;
        RECT 70.200 58.800 70.600 59.200 ;
        RECT 61.400 56.800 61.800 57.200 ;
        RECT 63.000 56.800 63.400 57.200 ;
        RECT 66.200 56.800 66.600 57.200 ;
        RECT 52.600 55.800 53.000 56.200 ;
        RECT 54.200 56.100 54.600 56.200 ;
        RECT 55.000 56.100 55.400 56.200 ;
        RECT 54.200 55.800 55.400 56.100 ;
        RECT 55.800 55.800 56.200 56.200 ;
        RECT 58.200 56.100 58.600 56.200 ;
        RECT 59.000 56.100 59.400 56.200 ;
        RECT 58.200 55.800 59.400 56.100 ;
        RECT 60.600 55.800 61.000 56.200 ;
        RECT 50.200 54.800 50.600 55.200 ;
        RECT 51.000 54.800 51.400 55.200 ;
        RECT 51.000 54.200 51.300 54.800 ;
        RECT 51.000 53.800 51.400 54.200 ;
        RECT 52.600 53.200 52.900 55.800 ;
        RECT 60.600 55.200 60.900 55.800 ;
        RECT 54.200 55.100 54.600 55.200 ;
        RECT 55.000 55.100 55.400 55.200 ;
        RECT 54.200 54.800 55.400 55.100 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 60.600 54.800 61.000 55.200 ;
        RECT 56.600 54.200 56.900 54.800 ;
        RECT 61.400 54.200 61.700 56.800 ;
        RECT 63.000 56.200 63.300 56.800 ;
        RECT 63.000 55.800 63.400 56.200 ;
        RECT 63.800 55.800 64.200 56.200 ;
        RECT 53.400 53.800 53.800 54.200 ;
        RECT 56.600 53.800 57.000 54.200 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 59.000 54.100 59.400 54.200 ;
        RECT 58.200 53.800 59.400 54.100 ;
        RECT 61.400 54.100 61.800 54.200 ;
        RECT 62.200 54.100 62.600 54.200 ;
        RECT 61.400 53.800 62.600 54.100 ;
        RECT 52.600 52.800 53.000 53.200 ;
        RECT 53.400 49.200 53.700 53.800 ;
        RECT 63.000 53.200 63.300 55.800 ;
        RECT 63.800 55.200 64.100 55.800 ;
        RECT 66.200 55.200 66.500 56.800 ;
        RECT 63.800 54.800 64.200 55.200 ;
        RECT 65.400 54.800 65.800 55.200 ;
        RECT 66.200 54.800 66.600 55.200 ;
        RECT 68.600 54.800 69.000 55.200 ;
        RECT 70.200 55.100 70.600 55.200 ;
        RECT 71.000 55.100 71.300 72.800 ;
        RECT 73.400 71.200 73.700 74.800 ;
        RECT 73.400 70.800 73.800 71.200 ;
        RECT 73.400 67.800 73.800 68.200 ;
        RECT 73.400 67.200 73.700 67.800 ;
        RECT 73.400 66.800 73.800 67.200 ;
        RECT 71.800 65.800 72.200 66.200 ;
        RECT 72.600 65.800 73.000 66.200 ;
        RECT 71.800 64.200 72.100 65.800 ;
        RECT 71.800 63.800 72.200 64.200 ;
        RECT 71.800 56.200 72.100 63.800 ;
        RECT 72.600 61.200 72.900 65.800 ;
        RECT 72.600 60.800 73.000 61.200 ;
        RECT 74.200 57.200 74.500 74.800 ;
        RECT 83.800 74.200 84.100 75.800 ;
        RECT 85.400 75.200 85.700 75.800 ;
        RECT 86.200 75.200 86.500 87.800 ;
        RECT 87.000 86.800 87.400 87.200 ;
        RECT 91.000 87.100 91.400 87.200 ;
        RECT 91.800 87.100 92.200 87.200 ;
        RECT 91.000 86.800 92.200 87.100 ;
        RECT 87.000 81.200 87.300 86.800 ;
        RECT 89.400 85.800 89.800 86.200 ;
        RECT 89.400 85.200 89.700 85.800 ;
        RECT 89.400 84.800 89.800 85.200 ;
        RECT 89.400 84.200 89.700 84.800 ;
        RECT 89.400 83.800 89.800 84.200 ;
        RECT 88.600 82.800 89.000 83.200 ;
        RECT 88.600 82.200 88.900 82.800 ;
        RECT 88.600 81.800 89.000 82.200 ;
        RECT 87.000 80.800 87.400 81.200 ;
        RECT 85.400 74.800 85.800 75.200 ;
        RECT 86.200 74.800 86.600 75.200 ;
        RECT 85.400 74.200 85.700 74.800 ;
        RECT 86.200 74.200 86.500 74.800 ;
        RECT 87.000 74.200 87.300 80.800 ;
        RECT 91.800 76.800 92.200 77.200 ;
        RECT 91.800 76.200 92.100 76.800 ;
        RECT 91.800 75.800 92.200 76.200 ;
        RECT 91.800 75.200 92.100 75.800 ;
        RECT 93.400 75.200 93.700 94.800 ;
        RECT 94.200 93.800 94.600 94.200 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 99.000 93.800 99.400 94.200 ;
        RECT 100.600 94.100 101.000 94.200 ;
        RECT 101.400 94.100 101.800 94.200 ;
        RECT 100.600 93.800 101.800 94.100 ;
        RECT 94.200 93.200 94.500 93.800 ;
        RECT 94.200 92.800 94.600 93.200 ;
        RECT 96.600 89.200 96.900 93.800 ;
        RECT 97.400 90.800 97.800 91.200 ;
        RECT 96.600 88.800 97.000 89.200 ;
        RECT 96.600 88.200 96.900 88.800 ;
        RECT 96.600 87.800 97.000 88.200 ;
        RECT 97.400 87.200 97.700 90.800 ;
        RECT 99.000 87.200 99.300 93.800 ;
        RECT 94.200 87.100 94.600 87.200 ;
        RECT 95.000 87.100 95.400 87.200 ;
        RECT 94.200 86.800 95.400 87.100 ;
        RECT 95.800 86.800 96.200 87.200 ;
        RECT 97.400 87.100 97.800 87.200 ;
        RECT 98.200 87.100 98.600 87.200 ;
        RECT 97.400 86.800 98.600 87.100 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 101.400 86.800 101.800 87.200 ;
        RECT 95.800 86.200 96.100 86.800 ;
        RECT 95.000 85.800 95.400 86.200 ;
        RECT 95.800 85.800 96.200 86.200 ;
        RECT 97.400 85.800 97.800 86.200 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 94.200 84.800 94.600 85.200 ;
        RECT 94.200 83.200 94.500 84.800 ;
        RECT 94.200 82.800 94.600 83.200 ;
        RECT 95.000 81.200 95.300 85.800 ;
        RECT 95.800 82.100 96.200 82.200 ;
        RECT 96.600 82.100 97.000 82.200 ;
        RECT 95.800 81.800 97.000 82.100 ;
        RECT 95.000 80.800 95.400 81.200 ;
        RECT 96.600 79.800 97.000 80.200 ;
        RECT 95.800 75.800 96.200 76.200 ;
        RECT 95.800 75.200 96.100 75.800 ;
        RECT 96.600 75.200 96.900 79.800 ;
        RECT 89.400 74.800 89.800 75.200 ;
        RECT 91.800 74.800 92.200 75.200 ;
        RECT 92.600 75.100 93.000 75.200 ;
        RECT 93.400 75.100 93.800 75.200 ;
        RECT 92.600 74.800 93.800 75.100 ;
        RECT 95.800 74.800 96.200 75.200 ;
        RECT 96.600 74.800 97.000 75.200 ;
        RECT 89.400 74.200 89.700 74.800 ;
        RECT 91.800 74.200 92.100 74.800 ;
        RECT 79.000 74.100 79.400 74.200 ;
        RECT 79.800 74.100 80.200 74.200 ;
        RECT 79.000 73.800 80.200 74.100 ;
        RECT 83.800 73.800 84.200 74.200 ;
        RECT 85.400 73.800 85.800 74.200 ;
        RECT 86.200 73.800 86.600 74.200 ;
        RECT 87.000 73.800 87.400 74.200 ;
        RECT 88.600 73.800 89.000 74.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 91.800 73.800 92.200 74.200 ;
        RECT 75.800 71.800 76.200 72.200 ;
        RECT 85.400 71.800 85.800 72.200 ;
        RECT 74.200 56.800 74.600 57.200 ;
        RECT 71.800 55.800 72.200 56.200 ;
        RECT 74.200 55.800 74.600 56.200 ;
        RECT 70.200 54.800 71.300 55.100 ;
        RECT 74.200 55.200 74.500 55.800 ;
        RECT 74.200 54.800 74.600 55.200 ;
        RECT 63.000 52.800 63.400 53.200 ;
        RECT 63.800 52.200 64.100 54.800 ;
        RECT 65.400 54.200 65.700 54.800 ;
        RECT 68.600 54.200 68.900 54.800 ;
        RECT 65.400 53.800 65.800 54.200 ;
        RECT 68.600 53.800 69.000 54.200 ;
        RECT 69.400 53.800 69.800 54.200 ;
        RECT 72.600 54.100 73.000 54.200 ;
        RECT 71.800 53.800 73.000 54.100 ;
        RECT 74.200 54.100 74.600 54.200 ;
        RECT 75.000 54.100 75.400 54.200 ;
        RECT 74.200 53.800 75.400 54.100 ;
        RECT 75.800 54.100 76.100 71.800 ;
        RECT 82.200 70.800 82.600 71.200 ;
        RECT 77.400 67.800 77.800 68.200 ;
        RECT 77.400 67.200 77.700 67.800 ;
        RECT 82.200 67.200 82.500 70.800 ;
        RECT 84.600 69.800 85.000 70.200 ;
        RECT 83.800 67.800 84.200 68.200 ;
        RECT 77.400 66.800 77.800 67.200 ;
        RECT 79.000 67.100 79.400 67.200 ;
        RECT 79.800 67.100 80.200 67.200 ;
        RECT 79.000 66.800 80.200 67.100 ;
        RECT 82.200 66.800 82.600 67.200 ;
        RECT 76.600 65.800 77.000 66.200 ;
        RECT 77.400 65.800 77.800 66.200 ;
        RECT 79.000 66.100 79.400 66.200 ;
        RECT 79.800 66.100 80.200 66.200 ;
        RECT 79.000 65.800 80.200 66.100 ;
        RECT 76.600 65.200 76.900 65.800 ;
        RECT 77.400 65.200 77.700 65.800 ;
        RECT 76.600 64.800 77.000 65.200 ;
        RECT 77.400 64.800 77.800 65.200 ;
        RECT 79.000 64.800 79.400 65.200 ;
        RECT 80.600 65.100 81.000 65.200 ;
        RECT 81.400 65.100 81.800 65.200 ;
        RECT 80.600 64.800 81.800 65.100 ;
        RECT 79.000 64.200 79.300 64.800 ;
        RECT 79.000 63.800 79.400 64.200 ;
        RECT 79.800 64.100 80.200 64.200 ;
        RECT 80.600 64.100 81.000 64.200 ;
        RECT 79.800 63.800 81.000 64.100 ;
        RECT 79.800 62.800 80.200 63.200 ;
        RECT 77.400 61.800 77.800 62.200 ;
        RECT 77.400 55.200 77.700 61.800 ;
        RECT 79.800 57.200 80.100 62.800 ;
        RECT 79.800 56.800 80.200 57.200 ;
        RECT 77.400 54.800 77.800 55.200 ;
        RECT 77.400 54.200 77.700 54.800 ;
        RECT 82.200 54.200 82.500 66.800 ;
        RECT 83.800 55.200 84.100 67.800 ;
        RECT 84.600 55.200 84.900 69.800 ;
        RECT 85.400 68.200 85.700 71.800 ;
        RECT 87.000 69.200 87.300 73.800 ;
        RECT 87.800 71.800 88.200 72.200 ;
        RECT 87.000 68.800 87.400 69.200 ;
        RECT 85.400 67.800 85.800 68.200 ;
        RECT 85.400 65.800 85.800 66.200 ;
        RECT 83.800 54.800 84.200 55.200 ;
        RECT 84.600 54.800 85.000 55.200 ;
        RECT 76.600 54.100 77.000 54.200 ;
        RECT 75.800 53.800 77.000 54.100 ;
        RECT 77.400 53.800 77.800 54.200 ;
        RECT 82.200 53.800 82.600 54.200 ;
        RECT 83.800 53.800 84.200 54.200 ;
        RECT 66.200 52.800 66.600 53.200 ;
        RECT 58.200 51.800 58.600 52.200 ;
        RECT 60.600 51.800 61.000 52.200 ;
        RECT 63.000 51.800 63.400 52.200 ;
        RECT 63.800 51.800 64.200 52.200 ;
        RECT 64.600 51.800 65.000 52.200 ;
        RECT 58.200 51.200 58.500 51.800 ;
        RECT 58.200 50.800 58.600 51.200 ;
        RECT 44.600 48.800 45.000 49.200 ;
        RECT 47.800 48.800 48.200 49.200 ;
        RECT 53.400 48.800 53.800 49.200 ;
        RECT 44.600 48.200 44.900 48.800 ;
        RECT 34.200 48.100 34.600 48.200 ;
        RECT 35.000 48.100 35.400 48.200 ;
        RECT 34.200 47.800 35.400 48.100 ;
        RECT 35.800 47.800 36.200 48.200 ;
        RECT 39.800 47.800 40.200 48.200 ;
        RECT 43.000 47.800 43.400 48.200 ;
        RECT 43.800 47.800 44.200 48.200 ;
        RECT 44.600 47.800 45.000 48.200 ;
        RECT 46.200 47.800 46.600 48.200 ;
        RECT 39.800 47.200 40.100 47.800 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 42.200 46.800 42.600 47.200 ;
        RECT 44.600 46.800 45.000 47.200 ;
        RECT 42.200 46.200 42.500 46.800 ;
        RECT 27.000 46.100 27.400 46.200 ;
        RECT 27.800 46.100 28.200 46.200 ;
        RECT 27.000 45.800 28.200 46.100 ;
        RECT 31.800 45.800 32.200 46.200 ;
        RECT 34.200 46.100 34.600 46.200 ;
        RECT 35.000 46.100 35.400 46.200 ;
        RECT 34.200 45.800 35.400 46.100 ;
        RECT 37.400 46.100 37.800 46.200 ;
        RECT 38.200 46.100 38.600 46.200 ;
        RECT 37.400 45.800 38.600 46.100 ;
        RECT 39.000 46.100 39.400 46.200 ;
        RECT 39.800 46.100 40.200 46.200 ;
        RECT 39.000 45.800 40.200 46.100 ;
        RECT 40.600 45.800 41.000 46.200 ;
        RECT 42.200 45.800 42.600 46.200 ;
        RECT 20.600 38.800 21.000 39.200 ;
        RECT 22.200 38.800 22.600 39.200 ;
        RECT 27.000 39.100 27.400 39.200 ;
        RECT 27.800 39.100 28.200 39.200 ;
        RECT 27.000 38.800 28.200 39.100 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 18.200 34.200 18.500 34.800 ;
        RECT 18.200 33.800 18.600 34.200 ;
        RECT 14.200 33.100 14.600 33.500 ;
        RECT 14.900 33.200 17.700 33.500 ;
        RECT 17.300 33.100 17.700 33.200 ;
        RECT 19.000 33.100 19.400 35.900 ;
        RECT 10.200 31.800 10.600 32.200 ;
        RECT 20.600 32.100 21.000 37.900 ;
        RECT 21.400 35.800 21.800 36.200 ;
        RECT 21.400 35.100 21.700 35.800 ;
        RECT 21.400 34.700 21.800 35.100 ;
        RECT 21.400 32.800 21.800 33.200 ;
        RECT 8.600 27.500 9.000 27.900 ;
        RECT 10.200 27.800 10.500 31.800 ;
        RECT 9.300 27.500 11.400 27.800 ;
        RECT 11.900 27.500 12.300 27.900 ;
        RECT 3.800 26.800 4.200 27.200 ;
        RECT 7.000 27.100 7.400 27.200 ;
        RECT 7.800 27.100 8.200 27.200 ;
        RECT 7.000 26.800 8.200 27.100 ;
        RECT 8.600 27.100 8.900 27.500 ;
        RECT 9.300 27.400 9.700 27.500 ;
        RECT 11.000 27.400 11.400 27.500 ;
        RECT 8.600 26.800 11.000 27.100 ;
        RECT 0.600 13.100 1.000 15.900 ;
        RECT 2.200 12.100 2.600 17.900 ;
        RECT 3.800 9.200 4.100 26.800 ;
        RECT 8.600 25.100 8.900 26.800 ;
        RECT 10.600 26.700 11.000 26.800 ;
        RECT 9.400 25.800 9.800 26.200 ;
        RECT 9.400 25.200 9.700 25.800 ;
        RECT 8.600 24.700 9.000 25.100 ;
        RECT 9.400 24.800 9.800 25.200 ;
        RECT 12.000 25.100 12.300 27.500 ;
        RECT 13.400 25.100 13.800 27.900 ;
        RECT 14.200 26.800 14.600 27.200 ;
        RECT 11.900 24.700 12.300 25.100 ;
        RECT 14.200 24.200 14.500 26.800 ;
        RECT 6.200 23.800 6.600 24.200 ;
        RECT 14.200 23.800 14.600 24.200 ;
        RECT 6.200 22.200 6.500 23.800 ;
        RECT 8.600 22.800 9.000 23.200 ;
        RECT 15.000 23.100 15.400 28.900 ;
        RECT 15.800 25.900 16.200 26.300 ;
        RECT 15.800 25.200 16.100 25.900 ;
        RECT 15.800 24.800 16.200 25.200 ;
        RECT 19.800 23.100 20.200 28.900 ;
        RECT 21.400 27.200 21.700 32.800 ;
        RECT 22.200 29.200 22.500 38.800 ;
        RECT 25.400 32.100 25.800 37.900 ;
        RECT 28.600 33.100 29.000 35.900 ;
        RECT 30.200 32.100 30.600 37.900 ;
        RECT 31.000 32.800 31.400 33.200 ;
        RECT 22.200 28.800 22.600 29.200 ;
        RECT 20.600 26.800 21.000 27.200 ;
        RECT 21.400 26.800 21.800 27.200 ;
        RECT 20.600 24.200 20.900 26.800 ;
        RECT 23.000 25.100 23.400 27.900 ;
        RECT 23.800 26.800 24.200 27.200 ;
        RECT 23.800 26.200 24.100 26.800 ;
        RECT 23.800 25.800 24.200 26.200 ;
        RECT 20.600 23.800 21.000 24.200 ;
        RECT 6.200 21.800 6.600 22.200 ;
        RECT 6.200 15.200 6.500 21.800 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 7.000 12.100 7.400 17.900 ;
        RECT 8.600 9.200 8.900 22.800 ;
        RECT 9.400 21.800 9.800 22.200 ;
        RECT 9.400 19.200 9.700 21.800 ;
        RECT 9.400 18.800 9.800 19.200 ;
        RECT 12.500 15.900 12.900 16.300 ;
        RECT 15.800 15.900 16.200 16.300 ;
        RECT 12.500 13.500 12.800 15.900 ;
        RECT 13.800 14.200 14.200 14.300 ;
        RECT 15.900 14.200 16.200 15.900 ;
        RECT 13.800 13.900 16.200 14.200 ;
        RECT 15.900 13.500 16.200 13.900 ;
        RECT 12.500 13.100 12.900 13.500 ;
        RECT 15.800 13.100 16.200 13.500 ;
        RECT 17.400 13.100 17.800 15.900 ;
        RECT 11.000 11.800 11.400 12.200 ;
        RECT 11.800 11.800 12.200 12.200 ;
        RECT 13.400 12.100 13.800 12.200 ;
        RECT 14.200 12.100 14.600 12.200 ;
        RECT 13.400 11.800 14.600 12.100 ;
        RECT 15.000 11.800 15.400 12.200 ;
        RECT 19.000 12.100 19.400 17.900 ;
        RECT 20.600 14.200 20.900 23.800 ;
        RECT 24.600 23.100 25.000 28.900 ;
        RECT 25.400 25.900 25.800 26.300 ;
        RECT 20.600 13.800 21.000 14.200 ;
        RECT 23.800 12.100 24.200 17.900 ;
        RECT 25.400 12.200 25.700 25.900 ;
        RECT 26.200 23.800 26.600 24.200 ;
        RECT 26.200 19.200 26.500 23.800 ;
        RECT 29.400 23.100 29.800 28.900 ;
        RECT 31.000 27.200 31.300 32.800 ;
        RECT 31.800 29.200 32.100 45.800 ;
        RECT 40.600 45.200 40.900 45.800 ;
        RECT 38.200 44.800 38.600 45.200 ;
        RECT 40.600 44.800 41.000 45.200 ;
        RECT 42.200 45.100 42.600 45.200 ;
        RECT 43.000 45.100 43.400 45.200 ;
        RECT 42.200 44.800 43.400 45.100 ;
        RECT 38.200 39.200 38.500 44.800 ;
        RECT 38.200 38.800 38.600 39.200 ;
        RECT 35.000 32.100 35.400 37.900 ;
        RECT 37.400 35.800 37.800 36.200 ;
        RECT 40.600 35.900 41.000 36.300 ;
        RECT 42.200 36.100 42.600 36.200 ;
        RECT 43.000 36.100 43.400 36.200 ;
        RECT 37.400 35.200 37.700 35.800 ;
        RECT 37.400 34.800 37.800 35.200 ;
        RECT 40.600 34.200 40.900 35.900 ;
        RECT 42.200 35.800 43.400 36.100 ;
        RECT 43.700 35.900 44.100 36.300 ;
        RECT 43.100 34.900 43.500 35.300 ;
        RECT 43.100 34.200 43.400 34.900 ;
        RECT 39.800 33.800 40.200 34.200 ;
        RECT 40.600 33.900 43.400 34.200 ;
        RECT 39.800 29.200 40.100 33.800 ;
        RECT 40.600 33.500 40.900 33.900 ;
        RECT 41.300 33.500 41.700 33.600 ;
        RECT 43.000 33.500 43.400 33.600 ;
        RECT 43.800 33.500 44.100 35.900 ;
        RECT 44.600 34.200 44.900 46.800 ;
        RECT 46.200 46.200 46.500 47.800 ;
        RECT 52.600 47.500 53.000 47.900 ;
        RECT 55.700 47.800 56.100 47.900 ;
        RECT 53.300 47.500 56.100 47.800 ;
        RECT 47.000 46.800 47.400 47.200 ;
        RECT 47.800 47.100 48.200 47.200 ;
        RECT 48.600 47.100 49.000 47.200 ;
        RECT 47.800 46.800 49.000 47.100 ;
        RECT 52.600 47.100 52.900 47.500 ;
        RECT 53.300 47.400 53.700 47.500 ;
        RECT 55.000 47.400 55.400 47.500 ;
        RECT 52.600 46.800 55.400 47.100 ;
        RECT 47.000 46.200 47.300 46.800 ;
        RECT 45.400 46.100 45.800 46.200 ;
        RECT 46.200 46.100 46.600 46.200 ;
        RECT 45.400 45.800 46.600 46.100 ;
        RECT 47.000 45.800 47.400 46.200 ;
        RECT 48.600 46.100 49.000 46.200 ;
        RECT 49.400 46.100 49.800 46.200 ;
        RECT 48.600 45.800 49.800 46.100 ;
        RECT 46.200 44.800 46.600 45.200 ;
        RECT 52.600 45.100 52.900 46.800 ;
        RECT 55.100 46.100 55.400 46.800 ;
        RECT 55.100 45.700 55.500 46.100 ;
        RECT 55.800 45.100 56.100 47.500 ;
        RECT 56.600 47.800 57.000 48.200 ;
        RECT 56.600 47.200 56.900 47.800 ;
        RECT 56.600 46.800 57.000 47.200 ;
        RECT 57.400 45.100 57.800 47.900 ;
        RECT 46.200 39.200 46.500 44.800 ;
        RECT 52.600 44.700 53.000 45.100 ;
        RECT 55.700 44.700 56.100 45.100 ;
        RECT 52.600 42.800 53.000 43.200 ;
        RECT 59.000 43.100 59.400 48.900 ;
        RECT 60.600 48.200 60.900 51.800 ;
        RECT 63.000 50.200 63.300 51.800 ;
        RECT 63.000 49.800 63.400 50.200 ;
        RECT 60.600 47.800 61.000 48.200 ;
        RECT 59.800 45.900 60.200 46.300 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 63.000 46.100 63.400 46.200 ;
        RECT 59.800 43.200 60.100 45.900 ;
        RECT 62.200 45.800 63.400 46.100 ;
        RECT 59.800 42.800 60.200 43.200 ;
        RECT 63.800 43.100 64.200 48.900 ;
        RECT 64.600 43.200 64.900 51.800 ;
        RECT 66.200 49.200 66.500 52.800 ;
        RECT 69.400 50.200 69.700 53.800 ;
        RECT 69.400 49.800 69.800 50.200 ;
        RECT 66.200 48.800 66.600 49.200 ;
        RECT 66.200 47.200 66.500 48.800 ;
        RECT 66.200 46.800 66.600 47.200 ;
        RECT 69.400 46.200 69.700 49.800 ;
        RECT 67.000 46.100 67.400 46.200 ;
        RECT 67.800 46.100 68.200 46.200 ;
        RECT 67.000 45.800 68.200 46.100 ;
        RECT 69.400 45.800 69.800 46.200 ;
        RECT 64.600 42.800 65.000 43.200 ;
        RECT 52.600 39.200 52.900 42.800 ;
        RECT 63.800 40.800 64.200 41.200 ;
        RECT 63.800 39.200 64.100 40.800 ;
        RECT 46.200 38.800 46.600 39.200 ;
        RECT 52.600 38.800 53.000 39.200 ;
        RECT 63.800 38.800 64.200 39.200 ;
        RECT 45.400 36.800 45.800 37.200 ;
        RECT 45.400 36.200 45.700 36.800 ;
        RECT 45.400 35.800 45.800 36.200 ;
        RECT 48.600 35.800 49.000 36.200 ;
        RECT 50.300 35.900 50.700 36.300 ;
        RECT 53.400 35.900 53.800 36.300 ;
        RECT 48.600 34.200 48.900 35.800 ;
        RECT 44.600 33.800 45.000 34.200 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 48.600 33.800 49.000 34.200 ;
        RECT 40.600 33.100 41.000 33.500 ;
        RECT 41.300 33.200 44.100 33.500 ;
        RECT 43.700 33.100 44.100 33.200 ;
        RECT 31.800 28.800 32.200 29.200 ;
        RECT 31.000 26.800 31.400 27.200 ;
        RECT 30.200 25.800 30.600 26.200 ;
        RECT 30.200 19.200 30.500 25.800 ;
        RECT 32.600 25.100 33.000 27.900 ;
        RECT 33.400 27.800 33.800 28.200 ;
        RECT 33.400 27.200 33.700 27.800 ;
        RECT 33.400 26.800 33.800 27.200 ;
        RECT 26.200 18.800 26.600 19.200 ;
        RECT 30.200 18.800 30.600 19.200 ;
        RECT 27.700 15.900 28.100 16.300 ;
        RECT 31.000 15.900 31.400 16.300 ;
        RECT 27.000 13.800 27.400 14.200 ;
        RECT 25.400 11.800 25.800 12.200 ;
        RECT 3.800 8.800 4.200 9.200 ;
        RECT 8.600 8.800 9.000 9.200 ;
        RECT 1.500 7.800 1.900 7.900 ;
        RECT 1.500 7.500 4.300 7.800 ;
        RECT 4.600 7.500 5.000 7.900 ;
        RECT 1.500 5.100 1.800 7.500 ;
        RECT 2.200 7.400 2.600 7.500 ;
        RECT 3.900 7.400 4.300 7.500 ;
        RECT 4.700 7.100 5.000 7.500 ;
        RECT 11.000 7.200 11.300 11.800 ;
        RECT 11.800 7.200 12.100 11.800 ;
        RECT 15.000 9.200 15.300 11.800 ;
        RECT 27.000 9.200 27.300 13.800 ;
        RECT 27.700 13.500 28.000 15.900 ;
        RECT 29.000 14.200 29.400 14.300 ;
        RECT 31.100 14.200 31.400 15.900 ;
        RECT 29.000 13.900 31.400 14.200 ;
        RECT 28.600 13.500 29.000 13.600 ;
        RECT 30.300 13.500 30.700 13.600 ;
        RECT 31.100 13.500 31.400 13.900 ;
        RECT 27.700 13.100 28.100 13.500 ;
        RECT 28.600 13.200 30.700 13.500 ;
        RECT 31.000 13.100 31.400 13.500 ;
        RECT 31.800 13.800 32.200 14.200 ;
        RECT 31.800 9.200 32.100 13.800 ;
        RECT 32.600 13.100 33.000 15.900 ;
        RECT 33.400 14.200 33.700 26.800 ;
        RECT 34.200 23.100 34.600 28.900 ;
        RECT 35.000 25.900 35.400 26.300 ;
        RECT 35.000 25.200 35.300 25.900 ;
        RECT 35.000 24.800 35.400 25.200 ;
        RECT 39.000 23.100 39.400 28.900 ;
        RECT 39.800 28.800 40.200 29.200 ;
        RECT 40.600 29.100 41.000 29.200 ;
        RECT 41.400 29.100 41.800 29.200 ;
        RECT 40.600 28.800 41.800 29.100 ;
        RECT 42.200 25.100 42.600 27.900 ;
        RECT 43.800 23.100 44.200 28.900 ;
        RECT 44.600 25.900 45.000 26.300 ;
        RECT 44.600 22.200 44.900 25.900 ;
        RECT 44.600 21.800 45.000 22.200 ;
        RECT 33.400 13.800 33.800 14.200 ;
        RECT 34.200 12.100 34.600 17.900 ;
        RECT 36.600 14.800 37.000 15.200 ;
        RECT 36.600 9.200 36.900 14.800 ;
        RECT 39.000 12.100 39.400 17.900 ;
        RECT 41.400 16.800 41.800 17.200 ;
        RECT 42.200 16.800 42.600 17.200 ;
        RECT 41.400 15.200 41.700 16.800 ;
        RECT 42.200 16.200 42.500 16.800 ;
        RECT 47.000 16.200 47.300 33.800 ;
        RECT 50.300 33.500 50.600 35.900 ;
        RECT 50.900 34.900 51.300 35.300 ;
        RECT 51.000 34.200 51.300 34.900 ;
        RECT 53.500 34.200 53.800 35.900 ;
        RECT 51.000 33.900 53.800 34.200 ;
        RECT 51.000 33.500 51.400 33.600 ;
        RECT 52.700 33.500 53.100 33.600 ;
        RECT 53.500 33.500 53.800 33.900 ;
        RECT 50.300 33.200 53.100 33.500 ;
        RECT 50.300 33.100 50.700 33.200 ;
        RECT 53.400 33.100 53.800 33.500 ;
        RECT 54.200 33.800 54.600 34.200 ;
        RECT 54.200 33.200 54.500 33.800 ;
        RECT 54.200 32.800 54.600 33.200 ;
        RECT 55.000 33.100 55.400 35.900 ;
        RECT 56.600 32.100 57.000 37.900 ;
        RECT 58.200 34.800 58.600 35.200 ;
        RECT 57.400 32.800 57.800 33.200 ;
        RECT 51.000 29.100 51.400 29.200 ;
        RECT 51.800 29.100 52.200 29.200 ;
        RECT 47.800 26.800 48.200 27.200 ;
        RECT 47.800 26.200 48.100 26.800 ;
        RECT 47.800 25.800 48.200 26.200 ;
        RECT 48.600 23.100 49.000 28.900 ;
        RECT 51.000 28.800 52.200 29.100 ;
        RECT 51.000 27.800 51.400 28.200 ;
        RECT 42.200 15.800 42.600 16.200 ;
        RECT 47.000 15.800 47.400 16.200 ;
        RECT 49.400 15.800 49.800 16.200 ;
        RECT 49.400 15.200 49.700 15.800 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 43.800 14.800 44.200 15.200 ;
        RECT 44.600 15.100 45.000 15.200 ;
        RECT 45.400 15.100 45.800 15.200 ;
        RECT 44.600 14.800 45.800 15.100 ;
        RECT 47.800 15.100 48.200 15.200 ;
        RECT 48.600 15.100 49.000 15.200 ;
        RECT 47.800 14.800 49.000 15.100 ;
        RECT 49.400 14.800 49.800 15.200 ;
        RECT 43.800 14.200 44.100 14.800 ;
        RECT 43.800 13.800 44.200 14.200 ;
        RECT 45.400 13.800 45.800 14.200 ;
        RECT 45.400 13.200 45.700 13.800 ;
        RECT 45.400 12.800 45.800 13.200 ;
        RECT 46.200 13.100 46.600 13.200 ;
        RECT 47.000 13.100 47.400 13.200 ;
        RECT 46.200 12.800 47.400 13.100 ;
        RECT 51.000 9.200 51.300 27.800 ;
        RECT 53.400 25.100 53.800 27.900 ;
        RECT 55.000 23.100 55.400 28.900 ;
        RECT 57.400 27.200 57.700 32.800 ;
        RECT 58.200 28.200 58.500 34.800 ;
        RECT 60.600 33.800 61.000 34.200 ;
        RECT 60.600 33.200 60.900 33.800 ;
        RECT 60.600 32.800 61.000 33.200 ;
        RECT 61.400 32.100 61.800 37.900 ;
        RECT 64.600 33.100 65.000 35.900 ;
        RECT 65.400 33.800 65.800 34.200 ;
        RECT 65.400 33.200 65.700 33.800 ;
        RECT 65.400 32.800 65.800 33.200 ;
        RECT 66.200 32.100 66.600 37.900 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 67.000 35.100 67.300 35.800 ;
        RECT 67.000 34.700 67.400 35.100 ;
        RECT 71.000 32.100 71.400 37.900 ;
        RECT 71.000 30.800 71.400 31.200 ;
        RECT 62.200 29.100 62.600 29.200 ;
        RECT 63.000 29.100 63.400 29.200 ;
        RECT 58.200 27.800 58.600 28.200 ;
        RECT 57.400 26.800 57.800 27.200 ;
        RECT 55.800 25.900 56.200 26.300 ;
        RECT 57.400 26.200 57.700 26.800 ;
        RECT 55.800 24.200 56.100 25.900 ;
        RECT 57.400 25.800 57.800 26.200 ;
        RECT 55.800 23.800 56.200 24.200 ;
        RECT 51.800 13.100 52.200 15.900 ;
        RECT 53.400 12.100 53.800 17.900 ;
        RECT 57.400 15.200 57.700 25.800 ;
        RECT 59.800 23.100 60.200 28.900 ;
        RECT 62.200 28.800 63.400 29.100 ;
        RECT 63.800 21.800 64.200 22.200 ;
        RECT 54.200 14.700 54.600 15.100 ;
        RECT 57.400 14.800 57.800 15.200 ;
        RECT 54.200 14.200 54.500 14.700 ;
        RECT 57.400 14.200 57.700 14.800 ;
        RECT 54.200 13.800 54.600 14.200 ;
        RECT 57.400 13.800 57.800 14.200 ;
        RECT 54.200 12.800 54.600 13.200 ;
        RECT 15.000 8.800 15.400 9.200 ;
        RECT 24.600 9.100 25.000 9.200 ;
        RECT 25.400 9.100 25.800 9.200 ;
        RECT 24.600 8.800 25.800 9.100 ;
        RECT 27.000 8.800 27.400 9.200 ;
        RECT 31.800 8.800 32.200 9.200 ;
        RECT 36.600 8.800 37.000 9.200 ;
        RECT 12.600 7.500 13.000 7.900 ;
        RECT 15.700 7.800 16.100 7.900 ;
        RECT 13.300 7.500 16.100 7.800 ;
        RECT 2.200 6.800 5.000 7.100 ;
        RECT 6.200 7.100 6.600 7.200 ;
        RECT 7.000 7.100 7.400 7.200 ;
        RECT 6.200 6.800 7.400 7.100 ;
        RECT 11.000 6.800 11.400 7.200 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 12.600 7.100 12.900 7.500 ;
        RECT 13.300 7.400 13.700 7.500 ;
        RECT 15.000 7.400 15.400 7.500 ;
        RECT 12.600 6.800 15.400 7.100 ;
        RECT 2.200 6.100 2.500 6.800 ;
        RECT 2.100 5.700 2.500 6.100 ;
        RECT 4.700 5.100 5.000 6.800 ;
        RECT 7.800 5.800 8.200 6.200 ;
        RECT 7.800 5.200 8.100 5.800 ;
        RECT 1.500 4.700 1.900 5.100 ;
        RECT 4.600 4.700 5.000 5.100 ;
        RECT 6.200 5.100 6.600 5.200 ;
        RECT 7.000 5.100 7.400 5.200 ;
        RECT 6.200 4.800 7.400 5.100 ;
        RECT 7.800 4.800 8.200 5.200 ;
        RECT 8.600 4.800 9.000 5.200 ;
        RECT 12.600 5.100 12.900 6.800 ;
        RECT 15.100 6.100 15.400 6.800 ;
        RECT 15.100 5.700 15.500 6.100 ;
        RECT 15.800 5.100 16.100 7.500 ;
        RECT 22.900 7.500 23.300 7.900 ;
        RECT 26.200 7.500 26.600 7.900 ;
        RECT 16.600 6.800 17.000 7.200 ;
        RECT 16.600 6.200 16.900 6.800 ;
        RECT 16.600 5.800 17.000 6.200 ;
        RECT 8.600 4.200 8.900 4.800 ;
        RECT 12.600 4.700 13.000 5.100 ;
        RECT 15.700 4.700 16.100 5.100 ;
        RECT 17.400 5.100 17.800 5.200 ;
        RECT 18.200 5.100 18.600 5.200 ;
        RECT 17.400 4.800 18.600 5.100 ;
        RECT 22.900 5.100 23.200 7.500 ;
        RECT 26.300 7.100 26.600 7.500 ;
        RECT 35.900 7.800 36.300 7.900 ;
        RECT 35.900 7.500 38.700 7.800 ;
        RECT 39.000 7.500 39.400 7.900 ;
        RECT 24.200 6.800 26.600 7.100 ;
        RECT 24.200 6.700 24.600 6.800 ;
        RECT 26.300 5.100 26.600 6.800 ;
        RECT 22.900 4.700 23.300 5.100 ;
        RECT 26.200 4.700 26.600 5.100 ;
        RECT 27.800 6.800 28.200 7.200 ;
        RECT 32.600 6.800 33.000 7.200 ;
        RECT 27.800 5.200 28.100 6.800 ;
        RECT 32.600 6.200 32.900 6.800 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 31.800 6.100 32.200 6.200 ;
        RECT 31.000 5.800 32.200 6.100 ;
        RECT 32.600 5.800 33.000 6.200 ;
        RECT 27.800 4.800 28.200 5.200 ;
        RECT 35.900 5.100 36.200 7.500 ;
        RECT 36.600 7.400 37.000 7.500 ;
        RECT 38.300 7.400 38.700 7.500 ;
        RECT 39.100 7.100 39.400 7.500 ;
        RECT 36.600 6.800 39.400 7.100 ;
        RECT 36.600 6.100 36.900 6.800 ;
        RECT 36.500 5.700 36.900 6.100 ;
        RECT 39.100 5.100 39.400 6.800 ;
        RECT 40.600 5.100 41.000 7.900 ;
        RECT 35.900 4.700 36.300 5.100 ;
        RECT 39.000 4.700 39.400 5.100 ;
        RECT 8.600 3.800 9.000 4.200 ;
        RECT 42.200 3.100 42.600 8.900 ;
        RECT 44.600 7.800 45.000 8.200 ;
        RECT 44.600 7.200 44.900 7.800 ;
        RECT 44.600 6.800 45.000 7.200 ;
        RECT 47.000 3.100 47.400 8.900 ;
        RECT 51.000 8.800 51.400 9.200 ;
        RECT 51.800 5.100 52.200 7.900 ;
        RECT 53.400 3.100 53.800 8.900 ;
        RECT 54.200 8.200 54.500 12.800 ;
        RECT 58.200 12.100 58.600 17.900 ;
        RECT 60.600 17.100 61.000 17.200 ;
        RECT 61.400 17.100 61.800 17.200 ;
        RECT 60.600 16.800 61.800 17.100 ;
        RECT 60.600 14.800 61.000 15.200 ;
        RECT 60.600 9.200 60.900 14.800 ;
        RECT 61.400 13.100 61.800 15.900 ;
        RECT 63.000 12.100 63.400 17.900 ;
        RECT 63.800 14.200 64.100 21.800 ;
        RECT 69.400 19.100 69.800 19.200 ;
        RECT 70.200 19.100 70.600 19.200 ;
        RECT 69.400 18.800 70.600 19.100 ;
        RECT 64.600 14.800 65.000 15.200 ;
        RECT 64.600 14.200 64.900 14.800 ;
        RECT 63.800 13.800 64.200 14.200 ;
        RECT 64.600 13.800 65.000 14.200 ;
        RECT 67.800 12.100 68.200 17.900 ;
        RECT 70.200 17.800 70.600 18.200 ;
        RECT 54.200 7.800 54.600 8.200 ;
        RECT 58.200 3.100 58.600 8.900 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 66.200 3.100 66.600 8.900 ;
        RECT 70.200 6.300 70.500 17.800 ;
        RECT 71.000 14.200 71.300 30.800 ;
        RECT 71.800 29.200 72.100 53.800 ;
        RECT 79.800 53.100 80.200 53.200 ;
        RECT 80.600 53.100 81.000 53.200 ;
        RECT 79.800 52.800 81.000 53.100 ;
        RECT 81.400 53.100 81.800 53.200 ;
        RECT 82.200 53.100 82.600 53.200 ;
        RECT 81.400 52.800 82.600 53.100 ;
        RECT 83.800 52.200 84.100 53.800 ;
        RECT 72.600 51.800 73.000 52.200 ;
        RECT 75.800 51.800 76.200 52.200 ;
        RECT 78.200 52.100 78.600 52.200 ;
        RECT 79.000 52.100 79.400 52.200 ;
        RECT 78.200 51.800 79.400 52.100 ;
        RECT 83.000 51.800 83.400 52.200 ;
        RECT 83.800 51.800 84.200 52.200 ;
        RECT 72.600 34.200 72.900 51.800 ;
        RECT 73.400 48.100 73.800 48.200 ;
        RECT 74.200 48.100 74.600 48.200 ;
        RECT 73.400 47.800 74.600 48.100 ;
        RECT 75.800 47.100 76.100 51.800 ;
        RECT 82.200 50.800 82.600 51.200 ;
        RECT 80.600 48.800 81.000 49.200 ;
        RECT 81.400 48.800 81.800 49.200 ;
        RECT 80.600 48.200 80.900 48.800 ;
        RECT 81.400 48.200 81.700 48.800 ;
        RECT 80.600 47.800 81.000 48.200 ;
        RECT 81.400 47.800 81.800 48.200 ;
        RECT 75.800 46.800 76.900 47.100 ;
        RECT 75.000 46.100 75.400 46.200 ;
        RECT 75.800 46.100 76.200 46.200 ;
        RECT 75.000 45.800 76.200 46.100 ;
        RECT 75.000 44.100 75.400 44.200 ;
        RECT 75.800 44.100 76.200 44.200 ;
        RECT 75.000 43.800 76.200 44.100 ;
        RECT 76.600 36.200 76.900 46.800 ;
        RECT 77.400 46.100 77.800 46.200 ;
        RECT 78.200 46.100 78.600 46.200 ;
        RECT 77.400 45.800 78.600 46.100 ;
        RECT 82.200 46.100 82.500 50.800 ;
        RECT 83.000 50.200 83.300 51.800 ;
        RECT 83.000 49.800 83.400 50.200 ;
        RECT 84.600 47.800 85.000 48.200 ;
        RECT 84.600 47.200 84.900 47.800 ;
        RECT 83.800 46.800 84.200 47.200 ;
        RECT 84.600 46.800 85.000 47.200 ;
        RECT 83.000 46.100 83.400 46.200 ;
        RECT 82.200 45.800 83.400 46.100 ;
        RECT 78.200 45.100 78.600 45.200 ;
        RECT 79.000 45.100 79.400 45.200 ;
        RECT 78.200 44.800 79.400 45.100 ;
        RECT 80.600 45.100 81.000 45.200 ;
        RECT 81.400 45.100 81.800 45.200 ;
        RECT 80.600 44.800 81.800 45.100 ;
        RECT 82.200 44.800 82.600 45.200 ;
        RECT 79.800 41.800 80.200 42.200 ;
        RECT 79.800 39.200 80.100 41.800 ;
        RECT 79.800 38.800 80.200 39.200 ;
        RECT 81.400 37.800 81.800 38.200 ;
        RECT 75.000 35.800 75.400 36.200 ;
        RECT 76.600 35.800 77.000 36.200 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 72.600 33.800 73.000 34.200 ;
        RECT 73.400 34.100 73.800 34.200 ;
        RECT 74.200 34.100 74.600 34.200 ;
        RECT 73.400 33.800 74.600 34.100 ;
        RECT 71.800 28.800 72.200 29.200 ;
        RECT 72.600 17.200 72.900 33.800 ;
        RECT 73.400 32.100 73.800 32.200 ;
        RECT 74.200 32.100 74.600 32.200 ;
        RECT 73.400 31.800 74.600 32.100 ;
        RECT 72.600 16.800 73.000 17.200 ;
        RECT 72.600 16.200 72.900 16.800 ;
        RECT 72.600 15.800 73.000 16.200 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 73.400 14.200 73.700 14.800 ;
        RECT 75.000 14.200 75.300 35.800 ;
        RECT 80.600 35.200 80.900 35.800 ;
        RECT 81.400 35.200 81.700 37.800 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 80.600 34.800 81.000 35.200 ;
        RECT 81.400 34.800 81.800 35.200 ;
        RECT 76.600 34.200 76.900 34.800 ;
        RECT 80.600 34.200 80.900 34.800 ;
        RECT 76.600 33.800 77.000 34.200 ;
        RECT 80.600 33.800 81.000 34.200 ;
        RECT 76.600 32.800 77.000 33.200 ;
        RECT 77.400 33.100 77.800 33.200 ;
        RECT 78.200 33.100 78.600 33.200 ;
        RECT 77.400 32.800 78.600 33.100 ;
        RECT 79.000 32.800 79.400 33.200 ;
        RECT 75.800 21.800 76.200 22.200 ;
        RECT 71.000 13.800 71.400 14.200 ;
        RECT 73.400 13.800 73.800 14.200 ;
        RECT 75.000 13.800 75.400 14.200 ;
        RECT 75.000 13.200 75.300 13.800 ;
        RECT 75.000 12.800 75.400 13.200 ;
        RECT 70.200 5.900 70.600 6.300 ;
        RECT 71.000 3.100 71.400 8.900 ;
        RECT 71.800 7.800 72.200 8.200 ;
        RECT 71.800 7.200 72.100 7.800 ;
        RECT 71.800 6.800 72.200 7.200 ;
        RECT 72.600 5.100 73.000 7.900 ;
        RECT 75.800 7.200 76.100 21.800 ;
        RECT 76.600 18.200 76.900 32.800 ;
        RECT 79.000 32.200 79.300 32.800 ;
        RECT 79.000 31.800 79.400 32.200 ;
        RECT 77.400 27.800 77.800 28.200 ;
        RECT 77.400 27.200 77.700 27.800 ;
        RECT 78.100 27.500 78.500 27.900 ;
        RECT 79.000 27.500 81.100 27.800 ;
        RECT 81.400 27.500 81.800 27.900 ;
        RECT 77.400 26.800 77.800 27.200 ;
        RECT 78.100 25.100 78.400 27.500 ;
        RECT 79.000 27.400 79.400 27.500 ;
        RECT 80.700 27.400 81.100 27.500 ;
        RECT 81.500 27.100 81.800 27.500 ;
        RECT 79.400 26.800 81.800 27.100 ;
        RECT 79.400 26.700 79.800 26.800 ;
        RECT 81.500 25.100 81.800 26.800 ;
        RECT 78.100 24.700 78.500 25.100 ;
        RECT 81.400 24.700 81.800 25.100 ;
        RECT 79.800 21.800 80.200 22.200 ;
        RECT 76.600 17.800 77.000 18.200 ;
        RECT 76.600 16.800 77.000 17.200 ;
        RECT 76.600 16.200 76.900 16.800 ;
        RECT 79.800 16.200 80.100 21.800 ;
        RECT 82.200 19.200 82.500 44.800 ;
        RECT 83.800 43.200 84.100 46.800 ;
        RECT 85.400 45.200 85.700 65.800 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 87.000 54.200 87.300 54.800 ;
        RECT 87.800 54.200 88.100 71.800 ;
        RECT 88.600 65.200 88.900 73.800 ;
        RECT 90.200 73.200 90.500 73.800 ;
        RECT 90.200 72.800 90.600 73.200 ;
        RECT 91.000 73.100 91.400 73.200 ;
        RECT 91.800 73.100 92.200 73.200 ;
        RECT 91.000 72.800 92.200 73.100 ;
        RECT 91.000 70.200 91.300 72.800 ;
        RECT 94.200 71.800 94.600 72.200 ;
        RECT 91.000 69.800 91.400 70.200 ;
        RECT 93.400 68.800 93.800 69.200 ;
        RECT 93.400 68.200 93.700 68.800 ;
        RECT 91.000 67.800 91.400 68.200 ;
        RECT 93.400 67.800 93.800 68.200 ;
        RECT 91.000 67.200 91.300 67.800 ;
        RECT 94.200 67.200 94.500 71.800 ;
        RECT 89.400 67.100 89.800 67.200 ;
        RECT 90.200 67.100 90.600 67.200 ;
        RECT 89.400 66.800 90.600 67.100 ;
        RECT 91.000 66.800 91.400 67.200 ;
        RECT 91.800 66.800 92.200 67.200 ;
        RECT 94.200 66.800 94.600 67.200 ;
        RECT 91.800 66.200 92.100 66.800 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 93.400 65.800 93.800 66.200 ;
        RECT 95.800 65.800 96.200 66.200 ;
        RECT 90.200 65.200 90.500 65.800 ;
        RECT 93.400 65.200 93.700 65.800 ;
        RECT 88.600 64.800 89.000 65.200 ;
        RECT 90.200 64.800 90.600 65.200 ;
        RECT 93.400 65.100 93.800 65.200 ;
        RECT 95.000 65.100 95.400 65.200 ;
        RECT 93.400 64.800 95.400 65.100 ;
        RECT 88.600 63.200 88.900 64.800 ;
        RECT 88.600 62.800 89.000 63.200 ;
        RECT 91.000 58.800 91.400 59.200 ;
        RECT 92.600 58.800 93.000 59.200 ;
        RECT 90.200 56.800 90.600 57.200 ;
        RECT 90.200 54.200 90.500 56.800 ;
        RECT 91.000 55.200 91.300 58.800 ;
        RECT 91.800 55.800 92.200 56.200 ;
        RECT 91.000 54.800 91.400 55.200 ;
        RECT 87.000 53.800 87.400 54.200 ;
        RECT 87.800 53.800 88.200 54.200 ;
        RECT 90.200 53.800 90.600 54.200 ;
        RECT 91.800 53.200 92.100 55.800 ;
        RECT 92.600 55.200 92.900 58.800 ;
        RECT 95.800 57.200 96.100 65.800 ;
        RECT 96.600 62.200 96.900 74.800 ;
        RECT 97.400 74.200 97.700 85.800 ;
        RECT 98.200 76.200 98.500 85.800 ;
        RECT 99.000 79.200 99.300 86.800 ;
        RECT 101.400 85.200 101.700 86.800 ;
        RECT 102.200 86.200 102.500 104.800 ;
        RECT 103.000 104.100 103.400 104.200 ;
        RECT 103.800 104.100 104.200 104.200 ;
        RECT 103.000 103.800 104.200 104.100 ;
        RECT 104.600 103.800 105.000 104.200 ;
        RECT 103.800 102.200 104.100 103.800 ;
        RECT 104.600 103.200 104.900 103.800 ;
        RECT 104.600 102.800 105.000 103.200 ;
        RECT 103.800 101.800 104.200 102.200 ;
        RECT 105.400 101.200 105.700 104.800 ;
        RECT 108.600 104.200 108.900 104.800 ;
        RECT 111.000 104.200 111.300 104.800 ;
        RECT 106.200 104.100 106.600 104.200 ;
        RECT 107.000 104.100 107.400 104.200 ;
        RECT 106.200 103.800 107.400 104.100 ;
        RECT 108.600 103.800 109.000 104.200 ;
        RECT 111.000 103.800 111.400 104.200 ;
        RECT 105.400 100.800 105.800 101.200 ;
        RECT 108.600 98.200 108.900 103.800 ;
        RECT 110.200 103.100 110.600 103.200 ;
        RECT 111.000 103.100 111.400 103.200 ;
        RECT 110.200 102.800 111.400 103.100 ;
        RECT 111.800 99.200 112.100 104.800 ;
        RECT 115.000 104.200 115.300 104.800 ;
        RECT 115.000 103.800 115.400 104.200 ;
        RECT 112.600 101.800 113.000 102.200 ;
        RECT 111.800 98.800 112.200 99.200 ;
        RECT 112.600 98.200 112.900 101.800 ;
        RECT 103.000 97.800 103.400 98.200 ;
        RECT 108.600 97.800 109.000 98.200 ;
        RECT 112.600 97.800 113.000 98.200 ;
        RECT 103.000 95.200 103.300 97.800 ;
        RECT 108.600 97.100 109.000 97.200 ;
        RECT 109.400 97.100 109.800 97.200 ;
        RECT 108.600 96.800 109.800 97.100 ;
        RECT 111.800 97.100 112.200 97.200 ;
        RECT 112.600 97.100 113.000 97.200 ;
        RECT 111.800 96.800 113.000 97.100 ;
        RECT 105.400 95.800 105.800 96.200 ;
        RECT 110.200 95.800 110.600 96.200 ;
        RECT 111.000 95.800 111.400 96.200 ;
        RECT 111.800 95.800 112.200 96.200 ;
        RECT 103.000 94.800 103.400 95.200 ;
        RECT 104.600 94.800 105.000 95.200 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 103.800 93.800 104.200 94.200 ;
        RECT 103.000 89.200 103.300 93.800 ;
        RECT 103.800 93.200 104.100 93.800 ;
        RECT 103.800 92.800 104.200 93.200 ;
        RECT 103.800 91.800 104.200 92.200 ;
        RECT 103.800 91.200 104.100 91.800 ;
        RECT 103.800 90.800 104.200 91.200 ;
        RECT 103.000 88.800 103.400 89.200 ;
        RECT 102.200 85.800 102.600 86.200 ;
        RECT 100.600 84.800 101.000 85.200 ;
        RECT 101.400 84.800 101.800 85.200 ;
        RECT 99.800 81.800 100.200 82.200 ;
        RECT 99.000 78.800 99.400 79.200 ;
        RECT 99.800 78.200 100.100 81.800 ;
        RECT 99.800 77.800 100.200 78.200 ;
        RECT 100.600 77.200 100.900 84.800 ;
        RECT 101.400 83.800 101.800 84.200 ;
        RECT 100.600 76.800 101.000 77.200 ;
        RECT 98.200 75.800 98.600 76.200 ;
        RECT 101.400 75.200 101.700 83.800 ;
        RECT 102.200 76.800 102.600 77.200 ;
        RECT 101.400 74.800 101.800 75.200 ;
        RECT 97.400 73.800 97.800 74.200 ;
        RECT 99.000 73.800 99.400 74.200 ;
        RECT 99.000 73.200 99.300 73.800 ;
        RECT 98.200 73.100 98.600 73.200 ;
        RECT 99.000 73.100 99.400 73.200 ;
        RECT 98.200 72.800 99.400 73.100 ;
        RECT 101.400 72.200 101.700 74.800 ;
        RECT 102.200 74.200 102.500 76.800 ;
        RECT 103.800 74.200 104.100 90.800 ;
        RECT 104.600 89.200 104.900 94.800 ;
        RECT 105.400 94.200 105.700 95.800 ;
        RECT 107.000 95.100 107.400 95.200 ;
        RECT 107.800 95.100 108.200 95.200 ;
        RECT 107.000 94.800 108.200 95.100 ;
        RECT 110.200 94.200 110.500 95.800 ;
        RECT 105.400 93.800 105.800 94.200 ;
        RECT 106.200 94.100 106.600 94.200 ;
        RECT 107.000 94.100 107.400 94.200 ;
        RECT 106.200 93.800 107.400 94.100 ;
        RECT 110.200 93.800 110.600 94.200 ;
        RECT 111.000 94.100 111.300 95.800 ;
        RECT 111.800 95.200 112.100 95.800 ;
        RECT 115.800 95.200 116.100 105.800 ;
        RECT 116.600 104.800 117.000 105.200 ;
        RECT 119.000 104.800 119.400 105.200 ;
        RECT 119.800 104.800 120.200 105.200 ;
        RECT 116.600 103.200 116.900 104.800 ;
        RECT 117.400 104.100 117.800 104.200 ;
        RECT 118.200 104.100 118.600 104.200 ;
        RECT 117.400 103.800 118.600 104.100 ;
        RECT 119.000 103.200 119.300 104.800 ;
        RECT 119.800 103.200 120.100 104.800 ;
        RECT 121.400 104.200 121.700 106.800 ;
        RECT 121.400 103.800 121.800 104.200 ;
        RECT 123.000 103.200 123.300 107.800 ;
        RECT 125.400 107.200 125.700 112.800 ;
        RECT 130.200 112.200 130.500 113.800 ;
        RECT 131.000 113.500 131.300 113.900 ;
        RECT 131.700 113.500 132.100 113.600 ;
        RECT 133.400 113.500 133.800 113.600 ;
        RECT 134.200 113.500 134.500 115.900 ;
        RECT 135.000 115.200 135.300 119.800 ;
        RECT 135.800 117.800 136.200 118.200 ;
        RECT 135.800 117.200 136.100 117.800 ;
        RECT 136.600 117.200 136.900 120.800 ;
        RECT 135.800 116.800 136.200 117.200 ;
        RECT 136.600 116.800 137.000 117.200 ;
        RECT 137.400 115.200 137.700 121.800 ;
        RECT 138.200 116.200 138.500 123.800 ;
        RECT 139.800 122.200 140.100 125.800 ;
        RECT 139.800 121.800 140.200 122.200 ;
        RECT 139.800 120.800 140.200 121.200 ;
        RECT 138.200 116.100 138.600 116.200 ;
        RECT 139.000 116.100 139.400 116.200 ;
        RECT 138.200 115.800 139.400 116.100 ;
        RECT 135.000 114.800 135.400 115.200 ;
        RECT 137.400 114.800 137.800 115.200 ;
        RECT 138.200 115.100 138.600 115.200 ;
        RECT 139.000 115.100 139.400 115.200 ;
        RECT 138.200 114.800 139.400 115.100 ;
        RECT 135.000 114.200 135.300 114.800 ;
        RECT 139.800 114.200 140.100 120.800 ;
        RECT 141.400 120.200 141.700 126.800 ;
        RECT 142.200 125.100 142.500 126.800 ;
        RECT 144.700 126.100 145.000 126.800 ;
        RECT 144.700 125.700 145.100 126.100 ;
        RECT 145.400 125.100 145.700 127.500 ;
        RECT 142.200 124.700 142.600 125.100 ;
        RECT 145.300 124.700 145.700 125.100 ;
        RECT 146.200 126.800 146.600 127.200 ;
        RECT 141.400 119.800 141.800 120.200 ;
        RECT 145.400 118.800 145.800 119.200 ;
        RECT 143.800 117.800 144.200 118.200 ;
        RECT 143.800 117.200 144.100 117.800 ;
        RECT 142.200 117.100 142.600 117.200 ;
        RECT 143.000 117.100 143.400 117.200 ;
        RECT 142.200 116.800 143.400 117.100 ;
        RECT 143.800 116.800 144.200 117.200 ;
        RECT 141.400 115.800 141.800 116.200 ;
        RECT 135.000 113.800 135.400 114.200 ;
        RECT 139.800 113.800 140.200 114.200 ;
        RECT 131.000 113.100 131.400 113.500 ;
        RECT 131.700 113.200 134.500 113.500 ;
        RECT 134.100 113.100 134.500 113.200 ;
        RECT 141.400 113.200 141.700 115.800 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 143.800 114.200 144.100 114.800 ;
        RECT 143.800 113.800 144.200 114.200 ;
        RECT 141.400 112.800 141.800 113.200 ;
        RECT 141.400 112.200 141.700 112.800 ;
        RECT 128.600 111.800 129.000 112.200 ;
        RECT 130.200 111.800 130.600 112.200 ;
        RECT 133.400 111.800 133.800 112.200 ;
        RECT 134.200 111.800 134.600 112.200 ;
        RECT 140.600 111.800 141.000 112.200 ;
        RECT 141.400 111.800 141.800 112.200 ;
        RECT 144.600 111.800 145.000 112.200 ;
        RECT 128.600 107.200 128.900 111.800 ;
        RECT 133.400 108.200 133.700 111.800 ;
        RECT 134.200 109.200 134.500 111.800 ;
        RECT 140.600 109.200 140.900 111.800 ;
        RECT 134.200 108.800 134.600 109.200 ;
        RECT 136.600 108.800 137.000 109.200 ;
        RECT 140.600 108.800 141.000 109.200 ;
        RECT 142.200 108.800 142.600 109.200 ;
        RECT 132.600 107.800 133.000 108.200 ;
        RECT 133.400 107.800 133.800 108.200 ;
        RECT 125.400 106.800 125.800 107.200 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 131.000 106.800 131.400 107.200 ;
        RECT 124.600 105.800 125.000 106.200 ;
        RECT 127.800 106.100 128.200 106.200 ;
        RECT 128.600 106.100 129.000 106.200 ;
        RECT 127.800 105.800 129.000 106.100 ;
        RECT 129.400 105.800 129.800 106.200 ;
        RECT 130.200 105.800 130.600 106.200 ;
        RECT 124.600 103.200 124.900 105.800 ;
        RECT 129.400 105.200 129.700 105.800 ;
        RECT 125.400 105.100 125.800 105.200 ;
        RECT 126.200 105.100 126.600 105.200 ;
        RECT 125.400 104.800 126.600 105.100 ;
        RECT 129.400 104.800 129.800 105.200 ;
        RECT 127.000 104.100 127.400 104.200 ;
        RECT 127.800 104.100 128.200 104.200 ;
        RECT 127.000 103.800 128.200 104.100 ;
        RECT 116.600 102.800 117.000 103.200 ;
        RECT 119.000 102.800 119.400 103.200 ;
        RECT 119.800 102.800 120.200 103.200 ;
        RECT 123.000 102.800 123.400 103.200 ;
        RECT 124.600 102.800 125.000 103.200 ;
        RECT 116.600 96.200 116.900 102.800 ;
        RECT 117.400 101.800 117.800 102.200 ;
        RECT 116.600 95.800 117.000 96.200 ;
        RECT 117.400 95.200 117.700 101.800 ;
        RECT 119.000 96.800 119.400 97.200 ;
        RECT 111.800 94.800 112.200 95.200 ;
        RECT 114.200 94.800 114.600 95.200 ;
        RECT 115.000 94.800 115.400 95.200 ;
        RECT 115.800 94.800 116.200 95.200 ;
        RECT 117.400 94.800 117.800 95.200 ;
        RECT 111.000 93.800 112.100 94.100 ;
        RECT 106.200 93.100 106.600 93.200 ;
        RECT 107.000 93.100 107.400 93.200 ;
        RECT 106.200 92.800 107.400 93.100 ;
        RECT 104.600 88.800 105.000 89.200 ;
        RECT 111.000 88.800 111.400 89.200 ;
        RECT 104.600 87.200 104.900 88.800 ;
        RECT 111.000 88.200 111.300 88.800 ;
        RECT 107.000 87.800 107.400 88.200 ;
        RECT 110.200 88.100 110.600 88.200 ;
        RECT 111.000 88.100 111.400 88.200 ;
        RECT 110.200 87.800 111.400 88.100 ;
        RECT 104.600 86.800 105.000 87.200 ;
        RECT 106.200 85.800 106.600 86.200 ;
        RECT 105.400 84.800 105.800 85.200 ;
        RECT 105.400 84.200 105.700 84.800 ;
        RECT 105.400 83.800 105.800 84.200 ;
        RECT 106.200 77.200 106.500 85.800 ;
        RECT 107.000 85.200 107.300 87.800 ;
        RECT 109.400 86.800 109.800 87.200 ;
        RECT 111.000 86.800 111.400 87.200 ;
        RECT 109.400 86.200 109.700 86.800 ;
        RECT 111.000 86.200 111.300 86.800 ;
        RECT 108.600 85.800 109.000 86.200 ;
        RECT 109.400 85.800 109.800 86.200 ;
        RECT 111.000 85.800 111.400 86.200 ;
        RECT 108.600 85.200 108.900 85.800 ;
        RECT 111.800 85.200 112.100 93.800 ;
        RECT 114.200 91.200 114.500 94.800 ;
        RECT 115.000 94.200 115.300 94.800 ;
        RECT 119.000 94.200 119.300 96.800 ;
        RECT 123.000 96.200 123.300 102.800 ;
        RECT 128.600 101.800 129.000 102.200 ;
        RECT 124.600 100.800 125.000 101.200 ;
        RECT 123.800 97.800 124.200 98.200 ;
        RECT 123.800 97.200 124.100 97.800 ;
        RECT 123.800 96.800 124.200 97.200 ;
        RECT 121.400 96.100 121.800 96.200 ;
        RECT 122.200 96.100 122.600 96.200 ;
        RECT 121.400 95.800 122.600 96.100 ;
        RECT 123.000 95.800 123.400 96.200 ;
        RECT 119.800 94.800 120.200 95.200 ;
        RECT 121.400 95.100 121.800 95.200 ;
        RECT 122.200 95.100 122.600 95.200 ;
        RECT 121.400 94.800 122.600 95.100 ;
        RECT 115.000 93.800 115.400 94.200 ;
        RECT 116.600 93.800 117.000 94.200 ;
        RECT 119.000 93.800 119.400 94.200 ;
        RECT 116.600 93.200 116.900 93.800 ;
        RECT 119.000 93.200 119.300 93.800 ;
        RECT 119.800 93.200 120.100 94.800 ;
        RECT 123.000 93.200 123.300 95.800 ;
        RECT 124.600 95.200 124.900 100.800 ;
        RECT 127.800 99.800 128.200 100.200 ;
        RECT 127.800 99.200 128.100 99.800 ;
        RECT 127.800 98.800 128.200 99.200 ;
        RECT 127.000 97.800 127.400 98.200 ;
        RECT 127.000 97.200 127.300 97.800 ;
        RECT 128.600 97.200 128.900 101.800 ;
        RECT 125.400 96.800 125.800 97.200 ;
        RECT 127.000 96.800 127.400 97.200 ;
        RECT 128.600 96.800 129.000 97.200 ;
        RECT 125.400 96.200 125.700 96.800 ;
        RECT 125.400 95.800 125.800 96.200 ;
        RECT 128.600 95.800 129.000 96.200 ;
        RECT 123.800 95.100 124.200 95.200 ;
        RECT 124.600 95.100 125.000 95.200 ;
        RECT 123.800 94.800 125.000 95.100 ;
        RECT 127.000 95.100 127.400 95.200 ;
        RECT 127.800 95.100 128.200 95.200 ;
        RECT 127.000 94.800 128.200 95.100 ;
        RECT 116.600 92.800 117.000 93.200 ;
        RECT 119.000 92.800 119.400 93.200 ;
        RECT 119.800 92.800 120.200 93.200 ;
        RECT 120.600 92.800 121.000 93.200 ;
        RECT 123.000 92.800 123.400 93.200 ;
        RECT 114.200 90.800 114.600 91.200 ;
        RECT 112.600 86.800 113.000 87.200 ;
        RECT 112.600 86.200 112.900 86.800 ;
        RECT 112.600 85.800 113.000 86.200 ;
        RECT 114.200 86.100 114.500 90.800 ;
        RECT 116.600 87.800 117.000 88.200 ;
        RECT 117.400 87.800 117.800 88.200 ;
        RECT 116.600 87.200 116.900 87.800 ;
        RECT 115.000 87.100 115.400 87.200 ;
        RECT 115.800 87.100 116.200 87.200 ;
        RECT 115.000 86.800 116.200 87.100 ;
        RECT 116.600 86.800 117.000 87.200 ;
        RECT 115.000 86.100 115.400 86.200 ;
        RECT 114.200 85.800 115.400 86.100 ;
        RECT 107.000 84.800 107.400 85.200 ;
        RECT 108.600 84.800 109.000 85.200 ;
        RECT 111.000 84.800 111.400 85.200 ;
        RECT 111.800 84.800 112.200 85.200 ;
        RECT 107.800 81.800 108.200 82.200 ;
        RECT 107.800 77.200 108.100 81.800 ;
        RECT 106.200 76.800 106.600 77.200 ;
        RECT 107.800 76.800 108.200 77.200 ;
        RECT 111.000 76.200 111.300 84.800 ;
        RECT 111.800 80.200 112.100 84.800 ;
        RECT 113.400 83.800 113.800 84.200 ;
        RECT 113.400 83.200 113.700 83.800 ;
        RECT 117.400 83.200 117.700 87.800 ;
        RECT 118.200 86.800 118.600 87.200 ;
        RECT 118.200 85.200 118.500 86.800 ;
        RECT 119.000 86.200 119.300 92.800 ;
        RECT 120.600 89.200 120.900 92.800 ;
        RECT 128.600 92.200 128.900 95.800 ;
        RECT 129.400 92.200 129.700 104.800 ;
        RECT 130.200 101.200 130.500 105.800 ;
        RECT 130.200 100.800 130.600 101.200 ;
        RECT 131.000 98.200 131.300 106.800 ;
        RECT 132.600 106.200 132.900 107.800 ;
        RECT 136.600 107.200 136.900 108.800 ;
        RECT 137.400 107.500 137.800 107.900 ;
        RECT 138.100 107.500 140.200 107.800 ;
        RECT 140.700 107.500 141.100 107.900 ;
        RECT 135.000 106.800 135.400 107.200 ;
        RECT 136.600 106.800 137.000 107.200 ;
        RECT 137.400 107.100 137.700 107.500 ;
        RECT 138.100 107.400 138.500 107.500 ;
        RECT 139.800 107.400 140.200 107.500 ;
        RECT 137.400 106.800 139.800 107.100 ;
        RECT 132.600 105.800 133.000 106.200 ;
        RECT 134.200 102.800 134.600 103.200 ;
        RECT 131.800 98.800 132.200 99.200 ;
        RECT 131.000 97.800 131.400 98.200 ;
        RECT 130.200 97.100 130.600 97.200 ;
        RECT 131.000 97.100 131.400 97.200 ;
        RECT 130.200 96.800 131.400 97.100 ;
        RECT 131.800 96.200 132.100 98.800 ;
        RECT 132.600 97.100 133.000 97.200 ;
        RECT 133.400 97.100 133.800 97.200 ;
        RECT 132.600 96.800 133.800 97.100 ;
        RECT 134.200 96.200 134.500 102.800 ;
        RECT 135.000 100.200 135.300 106.800 ;
        RECT 135.800 105.800 136.200 106.200 ;
        RECT 135.000 99.800 135.400 100.200 ;
        RECT 135.800 99.200 136.100 105.800 ;
        RECT 136.600 104.800 137.000 105.200 ;
        RECT 137.400 105.100 137.700 106.800 ;
        RECT 139.400 106.700 139.800 106.800 ;
        RECT 138.200 105.800 138.600 106.200 ;
        RECT 138.200 105.200 138.500 105.800 ;
        RECT 135.800 98.800 136.200 99.200 ;
        RECT 131.000 95.800 131.400 96.200 ;
        RECT 131.800 95.800 132.200 96.200 ;
        RECT 134.200 95.800 134.600 96.200 ;
        RECT 131.000 95.200 131.300 95.800 ;
        RECT 136.600 95.200 136.900 104.800 ;
        RECT 137.400 104.700 137.800 105.100 ;
        RECT 138.200 104.800 138.600 105.200 ;
        RECT 140.800 105.100 141.100 107.500 ;
        RECT 141.400 107.800 141.800 108.200 ;
        RECT 141.400 107.200 141.700 107.800 ;
        RECT 142.200 107.200 142.500 108.800 ;
        RECT 141.400 106.800 141.800 107.200 ;
        RECT 142.200 106.800 142.600 107.200 ;
        RECT 143.000 106.800 143.400 107.200 ;
        RECT 143.000 106.200 143.300 106.800 ;
        RECT 144.600 106.200 144.900 111.800 ;
        RECT 145.400 108.200 145.700 118.800 ;
        RECT 146.200 116.200 146.500 126.800 ;
        RECT 150.200 125.800 150.600 126.200 ;
        RECT 148.600 121.800 149.000 122.200 ;
        RECT 148.600 116.200 148.900 121.800 ;
        RECT 146.200 115.800 146.600 116.200 ;
        RECT 148.600 115.800 149.000 116.200 ;
        RECT 149.400 114.800 149.800 115.200 ;
        RECT 148.600 113.800 149.000 114.200 ;
        RECT 146.200 112.800 146.600 113.200 ;
        RECT 147.000 112.800 147.400 113.200 ;
        RECT 146.200 112.200 146.500 112.800 ;
        RECT 147.000 112.200 147.300 112.800 ;
        RECT 146.200 111.800 146.600 112.200 ;
        RECT 147.000 111.800 147.400 112.200 ;
        RECT 147.800 111.800 148.200 112.200 ;
        RECT 145.400 107.800 145.800 108.200 ;
        RECT 143.000 105.800 143.400 106.200 ;
        RECT 143.800 105.800 144.200 106.200 ;
        RECT 144.600 105.800 145.000 106.200 ;
        RECT 140.700 104.700 141.100 105.100 ;
        RECT 142.200 104.800 142.600 105.200 ;
        RECT 137.400 99.800 137.800 100.200 ;
        RECT 140.600 99.800 141.000 100.200 ;
        RECT 137.400 97.200 137.700 99.800 ;
        RECT 139.000 98.800 139.400 99.200 ;
        RECT 137.400 96.800 137.800 97.200 ;
        RECT 139.000 96.200 139.300 98.800 ;
        RECT 140.600 97.200 140.900 99.800 ;
        RECT 140.600 96.800 141.000 97.200 ;
        RECT 139.000 95.800 139.400 96.200 ;
        RECT 131.000 94.800 131.400 95.200 ;
        RECT 133.400 95.100 133.800 95.200 ;
        RECT 134.200 95.100 134.600 95.200 ;
        RECT 133.400 94.800 134.600 95.100 ;
        RECT 136.600 94.800 137.000 95.200 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 139.800 95.100 140.200 95.200 ;
        RECT 139.000 94.800 140.200 95.100 ;
        RECT 134.200 93.800 134.600 94.200 ;
        RECT 134.200 93.200 134.500 93.800 ;
        RECT 134.200 92.800 134.600 93.200 ;
        RECT 128.600 91.800 129.000 92.200 ;
        RECT 129.400 91.800 129.800 92.200 ;
        RECT 130.200 91.800 130.600 92.200 ;
        RECT 131.800 91.800 132.200 92.200 ;
        RECT 136.600 91.800 137.000 92.200 ;
        RECT 141.400 91.800 141.800 92.200 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 123.800 88.800 124.200 89.200 ;
        RECT 121.400 88.100 121.800 88.200 ;
        RECT 122.200 88.100 122.600 88.200 ;
        RECT 121.400 87.800 122.600 88.100 ;
        RECT 121.400 86.800 121.800 87.200 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 120.600 85.800 121.000 86.200 ;
        RECT 118.200 84.800 118.600 85.200 ;
        RECT 118.200 83.800 118.600 84.200 ;
        RECT 113.400 82.800 113.800 83.200 ;
        RECT 117.400 82.800 117.800 83.200 ;
        RECT 112.600 81.800 113.000 82.200 ;
        RECT 111.800 79.800 112.200 80.200 ;
        RECT 112.600 78.100 112.900 81.800 ;
        RECT 118.200 79.200 118.500 83.800 ;
        RECT 120.600 83.200 120.900 85.800 ;
        RECT 120.600 82.800 121.000 83.200 ;
        RECT 118.200 78.800 118.600 79.200 ;
        RECT 120.600 78.200 120.900 82.800 ;
        RECT 121.400 82.200 121.700 86.800 ;
        RECT 123.800 86.200 124.100 88.800 ;
        RECT 126.200 86.800 126.600 87.200 ;
        RECT 127.000 86.800 127.400 87.200 ;
        RECT 126.200 86.200 126.500 86.800 ;
        RECT 127.000 86.200 127.300 86.800 ;
        RECT 130.200 86.200 130.500 91.800 ;
        RECT 131.800 89.200 132.100 91.800 ;
        RECT 131.800 88.800 132.200 89.200 ;
        RECT 131.000 87.800 131.400 88.200 ;
        RECT 123.800 85.800 124.200 86.200 ;
        RECT 126.200 85.800 126.600 86.200 ;
        RECT 127.000 85.800 127.400 86.200 ;
        RECT 130.200 85.800 130.600 86.200 ;
        RECT 131.000 85.200 131.300 87.800 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 132.600 87.100 133.000 87.200 ;
        RECT 131.800 86.800 133.000 87.100 ;
        RECT 133.400 85.800 133.800 86.200 ;
        RECT 135.000 86.100 135.400 86.200 ;
        RECT 135.800 86.100 136.200 86.200 ;
        RECT 135.000 85.800 136.200 86.100 ;
        RECT 123.800 84.800 124.200 85.200 ;
        RECT 124.600 84.800 125.000 85.200 ;
        RECT 130.200 84.800 130.600 85.200 ;
        RECT 131.000 84.800 131.400 85.200 ;
        RECT 123.800 84.200 124.100 84.800 ;
        RECT 123.800 83.800 124.200 84.200 ;
        RECT 124.600 83.200 124.900 84.800 ;
        RECT 130.200 84.200 130.500 84.800 ;
        RECT 133.400 84.200 133.700 85.800 ;
        RECT 136.600 85.200 136.900 91.800 ;
        RECT 141.400 88.200 141.700 91.800 ;
        RECT 142.200 89.200 142.500 104.800 ;
        RECT 143.800 97.200 144.100 105.800 ;
        RECT 144.600 105.200 144.900 105.800 ;
        RECT 144.600 104.800 145.000 105.200 ;
        RECT 145.400 104.100 145.700 107.800 ;
        RECT 147.800 107.200 148.100 111.800 ;
        RECT 148.600 110.200 148.900 113.800 ;
        RECT 149.400 110.200 149.700 114.800 ;
        RECT 148.600 109.800 149.000 110.200 ;
        RECT 149.400 109.800 149.800 110.200 ;
        RECT 150.200 109.200 150.500 125.800 ;
        RECT 150.200 108.800 150.600 109.200 ;
        RECT 149.400 107.800 149.800 108.200 ;
        RECT 151.000 107.800 151.400 108.200 ;
        RECT 149.400 107.200 149.700 107.800 ;
        RECT 147.800 106.800 148.200 107.200 ;
        RECT 149.400 106.800 149.800 107.200 ;
        RECT 150.200 106.800 150.600 107.200 ;
        RECT 146.200 106.100 146.600 106.200 ;
        RECT 147.000 106.100 147.400 106.200 ;
        RECT 148.600 106.100 149.000 106.200 ;
        RECT 146.200 105.800 149.000 106.100 ;
        RECT 147.800 105.100 148.200 105.200 ;
        RECT 148.600 105.100 149.000 105.200 ;
        RECT 147.800 104.800 149.000 105.100 ;
        RECT 146.200 104.100 146.600 104.200 ;
        RECT 145.400 103.800 146.600 104.100 ;
        RECT 147.000 101.800 147.400 102.200 ;
        RECT 143.800 96.800 144.200 97.200 ;
        RECT 147.000 96.200 147.300 101.800 ;
        RECT 147.800 97.100 148.200 97.200 ;
        RECT 148.600 97.100 149.000 97.200 ;
        RECT 147.800 96.800 149.000 97.100 ;
        RECT 150.200 96.200 150.500 106.800 ;
        RECT 151.000 105.200 151.300 107.800 ;
        RECT 151.000 104.800 151.400 105.200 ;
        RECT 147.000 95.800 147.400 96.200 ;
        RECT 150.200 95.800 150.600 96.200 ;
        RECT 150.200 95.200 150.500 95.800 ;
        RECT 147.000 94.800 147.400 95.200 ;
        RECT 148.600 95.100 149.000 95.200 ;
        RECT 149.400 95.100 149.800 95.200 ;
        RECT 148.600 94.800 149.800 95.100 ;
        RECT 150.200 94.800 150.600 95.200 ;
        RECT 147.000 94.200 147.300 94.800 ;
        RECT 143.000 93.800 143.400 94.200 ;
        RECT 145.400 94.100 145.800 94.200 ;
        RECT 146.200 94.100 146.600 94.200 ;
        RECT 145.400 93.800 146.600 94.100 ;
        RECT 147.000 93.800 147.400 94.200 ;
        RECT 143.000 93.200 143.300 93.800 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 144.600 92.800 145.000 93.200 ;
        RECT 143.000 89.200 143.300 92.800 ;
        RECT 143.800 91.800 144.200 92.200 ;
        RECT 143.800 90.200 144.100 91.800 ;
        RECT 143.800 89.800 144.200 90.200 ;
        RECT 142.200 88.800 142.600 89.200 ;
        RECT 143.000 88.800 143.400 89.200 ;
        RECT 144.600 88.200 144.900 92.800 ;
        RECT 146.200 91.800 146.600 92.200 ;
        RECT 141.400 87.800 141.800 88.200 ;
        RECT 143.000 87.800 143.400 88.200 ;
        RECT 143.800 87.800 144.200 88.200 ;
        RECT 144.600 87.800 145.000 88.200 ;
        RECT 140.600 87.100 141.000 87.200 ;
        RECT 141.400 87.100 141.800 87.200 ;
        RECT 140.600 86.800 141.800 87.100 ;
        RECT 143.000 86.200 143.300 87.800 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 139.000 85.800 139.400 86.200 ;
        RECT 143.000 85.800 143.400 86.200 ;
        RECT 136.600 84.800 137.000 85.200 ;
        RECT 136.600 84.200 136.900 84.800 ;
        RECT 138.200 84.200 138.500 85.800 ;
        RECT 139.000 85.200 139.300 85.800 ;
        RECT 143.800 85.200 144.100 87.800 ;
        RECT 146.200 87.200 146.500 91.800 ;
        RECT 147.800 88.800 148.200 89.200 ;
        RECT 146.200 86.800 146.600 87.200 ;
        RECT 147.800 86.200 148.100 88.800 ;
        RECT 148.600 87.800 149.000 88.200 ;
        RECT 144.600 86.100 145.000 86.200 ;
        RECT 145.400 86.100 145.800 86.200 ;
        RECT 144.600 85.800 145.800 86.100 ;
        RECT 147.800 85.800 148.200 86.200 ;
        RECT 139.000 84.800 139.400 85.200 ;
        RECT 139.800 84.800 140.200 85.200 ;
        RECT 143.800 84.800 144.200 85.200 ;
        RECT 146.200 85.100 146.600 85.200 ;
        RECT 147.000 85.100 147.400 85.200 ;
        RECT 146.200 84.800 147.400 85.100 ;
        RECT 139.800 84.200 140.100 84.800 ;
        RECT 148.600 84.200 148.900 87.800 ;
        RECT 130.200 83.800 130.600 84.200 ;
        RECT 133.400 83.800 133.800 84.200 ;
        RECT 135.000 83.800 135.400 84.200 ;
        RECT 136.600 83.800 137.000 84.200 ;
        RECT 138.200 83.800 138.600 84.200 ;
        RECT 139.800 83.800 140.200 84.200 ;
        RECT 145.400 84.100 145.800 84.200 ;
        RECT 146.200 84.100 146.600 84.200 ;
        RECT 145.400 83.800 146.600 84.100 ;
        RECT 147.000 83.800 147.400 84.200 ;
        RECT 148.600 83.800 149.000 84.200 ;
        RECT 135.000 83.200 135.300 83.800 ;
        RECT 124.600 82.800 125.000 83.200 ;
        RECT 130.200 82.800 130.600 83.200 ;
        RECT 135.000 82.800 135.400 83.200 ;
        RECT 121.400 81.800 121.800 82.200 ;
        RECT 126.200 81.800 126.600 82.200 ;
        RECT 128.600 81.800 129.000 82.200 ;
        RECT 126.200 78.200 126.500 81.800 ;
        RECT 112.600 77.800 113.700 78.100 ;
        RECT 111.800 77.100 112.200 77.200 ;
        RECT 112.600 77.100 113.000 77.200 ;
        RECT 111.800 76.800 113.000 77.100 ;
        RECT 113.400 76.200 113.700 77.800 ;
        RECT 114.200 77.800 114.600 78.200 ;
        RECT 119.000 77.800 119.400 78.200 ;
        RECT 120.600 77.800 121.000 78.200 ;
        RECT 126.200 77.800 126.600 78.200 ;
        RECT 128.600 78.100 128.900 81.800 ;
        RECT 130.200 79.200 130.500 82.800 ;
        RECT 135.800 81.800 136.200 82.200 ;
        RECT 139.000 81.800 139.400 82.200 ;
        RECT 143.000 81.800 143.400 82.200 ;
        RECT 144.600 81.800 145.000 82.200 ;
        RECT 135.800 81.200 136.100 81.800 ;
        RECT 135.800 80.800 136.200 81.200 ;
        RECT 139.000 80.200 139.300 81.800 ;
        RECT 141.400 80.800 141.800 81.200 ;
        RECT 139.000 79.800 139.400 80.200 ;
        RECT 130.200 78.800 130.600 79.200 ;
        RECT 139.000 78.800 139.400 79.200 ;
        RECT 127.800 77.800 128.900 78.100 ;
        RECT 139.000 78.200 139.300 78.800 ;
        RECT 139.000 77.800 139.400 78.200 ;
        RECT 139.800 77.800 140.200 78.200 ;
        RECT 114.200 76.200 114.500 77.800 ;
        RECT 115.000 77.100 115.400 77.200 ;
        RECT 115.800 77.100 116.200 77.200 ;
        RECT 115.000 76.800 116.200 77.100 ;
        RECT 111.000 75.800 111.400 76.200 ;
        RECT 113.400 75.800 113.800 76.200 ;
        RECT 114.200 75.800 114.600 76.200 ;
        RECT 116.600 75.800 117.000 76.200 ;
        RECT 111.000 75.200 111.300 75.800 ;
        RECT 113.400 75.200 113.700 75.800 ;
        RECT 116.600 75.200 116.900 75.800 ;
        RECT 107.800 75.100 108.200 75.200 ;
        RECT 108.600 75.100 109.000 75.200 ;
        RECT 107.800 74.800 109.000 75.100 ;
        RECT 111.000 74.800 111.400 75.200 ;
        RECT 112.600 74.800 113.000 75.200 ;
        RECT 113.400 74.800 113.800 75.200 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 102.200 73.800 102.600 74.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 107.000 73.800 107.400 74.200 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 109.400 74.100 109.800 74.200 ;
        RECT 108.600 73.800 109.800 74.100 ;
        RECT 107.000 73.200 107.300 73.800 ;
        RECT 111.000 73.200 111.300 74.800 ;
        RECT 112.600 74.200 112.900 74.800 ;
        RECT 119.000 74.200 119.300 77.800 ;
        RECT 127.800 77.200 128.100 77.800 ;
        RECT 139.800 77.200 140.100 77.800 ;
        RECT 141.400 77.200 141.700 80.800 ;
        RECT 121.400 77.100 121.800 77.200 ;
        RECT 122.200 77.100 122.600 77.200 ;
        RECT 121.400 76.800 122.600 77.100 ;
        RECT 123.800 76.800 124.200 77.200 ;
        RECT 127.800 76.800 128.200 77.200 ;
        RECT 128.600 76.800 129.000 77.200 ;
        RECT 138.200 76.800 138.600 77.200 ;
        RECT 139.000 76.800 139.400 77.200 ;
        RECT 139.800 76.800 140.200 77.200 ;
        RECT 141.400 76.800 141.800 77.200 ;
        RECT 142.200 76.800 142.600 77.200 ;
        RECT 119.800 75.800 120.200 76.200 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 119.000 73.800 119.400 74.200 ;
        RECT 119.800 73.200 120.100 75.800 ;
        RECT 120.600 74.800 121.000 75.200 ;
        RECT 122.200 75.100 122.600 75.200 ;
        RECT 123.000 75.100 123.400 75.200 ;
        RECT 122.200 74.800 123.400 75.100 ;
        RECT 120.600 74.200 120.900 74.800 ;
        RECT 123.800 74.200 124.100 76.800 ;
        RECT 128.600 76.200 128.900 76.800 ;
        RECT 126.200 75.800 126.600 76.200 ;
        RECT 127.000 75.800 127.400 76.200 ;
        RECT 128.600 75.800 129.000 76.200 ;
        RECT 131.000 76.100 131.400 76.200 ;
        RECT 131.800 76.100 132.200 76.200 ;
        RECT 131.000 75.800 132.200 76.100 ;
        RECT 133.300 75.900 133.700 76.300 ;
        RECT 136.600 75.900 137.000 76.300 ;
        RECT 120.600 73.800 121.000 74.200 ;
        RECT 123.800 73.800 124.200 74.200 ;
        RECT 124.600 74.100 125.000 74.200 ;
        RECT 125.400 74.100 125.800 74.200 ;
        RECT 124.600 73.800 125.800 74.100 ;
        RECT 126.200 73.200 126.500 75.800 ;
        RECT 127.000 75.200 127.300 75.800 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 130.200 74.800 130.600 75.200 ;
        RECT 128.600 74.100 129.000 74.200 ;
        RECT 129.400 74.100 129.800 74.200 ;
        RECT 128.600 73.800 129.800 74.100 ;
        RECT 103.800 73.100 104.200 73.200 ;
        RECT 104.600 73.100 105.000 73.200 ;
        RECT 103.800 72.800 105.000 73.100 ;
        RECT 105.400 73.100 105.800 73.200 ;
        RECT 106.200 73.100 106.600 73.200 ;
        RECT 105.400 72.800 106.600 73.100 ;
        RECT 107.000 72.800 107.400 73.200 ;
        RECT 111.000 72.800 111.400 73.200 ;
        RECT 112.600 72.800 113.000 73.200 ;
        RECT 119.800 72.800 120.200 73.200 ;
        RECT 120.600 72.800 121.000 73.200 ;
        RECT 124.600 73.100 125.000 73.200 ;
        RECT 125.400 73.100 125.800 73.200 ;
        RECT 124.600 72.800 125.800 73.100 ;
        RECT 126.200 72.800 126.600 73.200 ;
        RECT 98.200 71.800 98.600 72.200 ;
        RECT 101.400 71.800 101.800 72.200 ;
        RECT 103.000 71.800 103.400 72.200 ;
        RECT 107.800 71.800 108.200 72.200 ;
        RECT 111.000 71.800 111.400 72.200 ;
        RECT 98.200 68.100 98.500 71.800 ;
        RECT 103.000 69.200 103.300 71.800 ;
        RECT 97.400 67.800 98.500 68.100 ;
        RECT 99.000 68.800 99.400 69.200 ;
        RECT 103.000 68.800 103.400 69.200 ;
        RECT 97.400 66.200 97.700 67.800 ;
        RECT 98.200 67.100 98.600 67.200 ;
        RECT 99.000 67.100 99.300 68.800 ;
        RECT 107.800 68.200 108.100 71.800 ;
        RECT 107.800 67.800 108.200 68.200 ;
        RECT 107.800 67.200 108.100 67.800 ;
        RECT 111.000 67.200 111.300 71.800 ;
        RECT 112.600 69.200 112.900 72.800 ;
        RECT 115.800 71.800 116.200 72.200 ;
        RECT 112.600 68.800 113.000 69.200 ;
        RECT 112.600 68.100 113.000 68.200 ;
        RECT 113.400 68.100 113.800 68.200 ;
        RECT 112.600 67.800 113.800 68.100 ;
        RECT 115.000 67.800 115.400 68.200 ;
        RECT 98.200 66.800 99.300 67.100 ;
        RECT 103.000 66.800 103.400 67.200 ;
        RECT 106.200 66.800 106.600 67.200 ;
        RECT 107.800 66.800 108.200 67.200 ;
        RECT 111.000 66.800 111.400 67.200 ;
        RECT 97.400 65.800 97.800 66.200 ;
        RECT 103.000 65.200 103.300 66.800 ;
        RECT 106.200 66.200 106.500 66.800 ;
        RECT 115.000 66.200 115.300 67.800 ;
        RECT 115.800 66.200 116.100 71.800 ;
        RECT 119.800 69.200 120.100 72.800 ;
        RECT 119.800 68.800 120.200 69.200 ;
        RECT 119.000 67.800 119.400 68.200 ;
        RECT 119.000 66.200 119.300 67.800 ;
        RECT 120.600 67.200 120.900 72.800 ;
        RECT 121.400 71.800 121.800 72.200 ;
        RECT 121.400 68.200 121.700 71.800 ;
        RECT 126.200 69.100 126.600 69.200 ;
        RECT 126.200 68.800 127.300 69.100 ;
        RECT 126.200 68.200 126.500 68.800 ;
        RECT 121.400 67.800 121.800 68.200 ;
        RECT 124.600 67.800 125.000 68.200 ;
        RECT 125.400 67.800 125.800 68.200 ;
        RECT 126.200 67.800 126.600 68.200 ;
        RECT 124.600 67.200 124.900 67.800 ;
        RECT 125.400 67.200 125.700 67.800 ;
        RECT 120.600 66.800 121.000 67.200 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 122.200 66.800 122.600 67.200 ;
        RECT 124.600 66.800 125.000 67.200 ;
        RECT 125.400 66.800 125.800 67.200 ;
        RECT 103.800 66.100 104.200 66.200 ;
        RECT 104.600 66.100 105.000 66.200 ;
        RECT 103.800 65.800 105.000 66.100 ;
        RECT 106.200 65.800 106.600 66.200 ;
        RECT 110.200 65.800 110.600 66.200 ;
        RECT 115.000 65.800 115.400 66.200 ;
        RECT 115.800 65.800 116.200 66.200 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 110.200 65.200 110.500 65.800 ;
        RECT 120.600 65.200 120.900 66.800 ;
        RECT 121.400 66.200 121.700 66.800 ;
        RECT 121.400 65.800 121.800 66.200 ;
        RECT 103.000 65.100 103.400 65.200 ;
        RECT 104.600 65.100 105.000 65.200 ;
        RECT 103.000 64.800 105.000 65.100 ;
        RECT 110.200 64.800 110.600 65.200 ;
        RECT 114.200 64.800 114.600 65.200 ;
        RECT 115.800 64.800 116.200 65.200 ;
        RECT 117.400 65.100 117.800 65.200 ;
        RECT 118.200 65.100 118.600 65.200 ;
        RECT 117.400 64.800 118.600 65.100 ;
        RECT 119.000 65.100 119.400 65.200 ;
        RECT 119.800 65.100 120.200 65.200 ;
        RECT 119.000 64.800 120.200 65.100 ;
        RECT 120.600 64.800 121.000 65.200 ;
        RECT 114.200 64.200 114.500 64.800 ;
        RECT 115.800 64.200 116.100 64.800 ;
        RECT 122.200 64.200 122.500 66.800 ;
        RECT 123.000 66.100 123.400 66.200 ;
        RECT 123.800 66.100 124.200 66.200 ;
        RECT 123.000 65.800 124.200 66.100 ;
        RECT 127.000 65.200 127.300 68.800 ;
        RECT 127.800 66.100 128.200 66.200 ;
        RECT 128.600 66.100 129.000 66.200 ;
        RECT 127.800 65.800 129.000 66.100 ;
        RECT 130.200 65.200 130.500 74.800 ;
        RECT 131.000 66.200 131.300 75.800 ;
        RECT 132.600 73.800 133.000 74.200 ;
        RECT 131.000 65.800 131.400 66.200 ;
        RECT 127.000 64.800 127.400 65.200 ;
        RECT 128.600 64.800 129.000 65.200 ;
        RECT 129.400 65.100 129.800 65.200 ;
        RECT 130.200 65.100 130.600 65.200 ;
        RECT 129.400 64.800 130.600 65.100 ;
        RECT 131.000 65.100 131.400 65.200 ;
        RECT 131.800 65.100 132.200 65.200 ;
        RECT 131.000 64.800 132.200 65.100 ;
        RECT 128.600 64.200 128.900 64.800 ;
        RECT 114.200 63.800 114.600 64.200 ;
        RECT 115.800 63.800 116.200 64.200 ;
        RECT 122.200 63.800 122.600 64.200 ;
        RECT 128.600 63.800 129.000 64.200 ;
        RECT 96.600 61.800 97.000 62.200 ;
        RECT 99.000 61.800 99.400 62.200 ;
        RECT 106.200 61.800 106.600 62.200 ;
        RECT 108.600 61.800 109.000 62.200 ;
        RECT 115.000 61.800 115.400 62.200 ;
        RECT 117.400 61.800 117.800 62.200 ;
        RECT 131.000 61.800 131.400 62.200 ;
        RECT 98.200 60.800 98.600 61.200 ;
        RECT 93.400 57.100 93.800 57.200 ;
        RECT 94.200 57.100 94.600 57.200 ;
        RECT 93.400 56.800 94.600 57.100 ;
        RECT 95.800 56.800 96.200 57.200 ;
        RECT 94.200 55.800 94.600 56.200 ;
        RECT 94.200 55.200 94.500 55.800 ;
        RECT 95.800 55.200 96.100 56.800 ;
        RECT 97.400 56.100 97.800 56.200 ;
        RECT 98.200 56.100 98.500 60.800 ;
        RECT 99.000 57.200 99.300 61.800 ;
        RECT 106.200 59.200 106.500 61.800 ;
        RECT 108.600 61.200 108.900 61.800 ;
        RECT 108.600 60.800 109.000 61.200 ;
        RECT 106.200 58.800 106.600 59.200 ;
        RECT 109.400 59.100 109.800 59.200 ;
        RECT 108.600 58.800 109.800 59.100 ;
        RECT 112.600 58.800 113.000 59.200 ;
        RECT 103.800 57.800 104.200 58.200 ;
        RECT 107.800 57.800 108.200 58.200 ;
        RECT 103.800 57.200 104.100 57.800 ;
        RECT 99.000 56.800 99.400 57.200 ;
        RECT 103.800 56.800 104.200 57.200 ;
        RECT 106.200 57.100 106.600 57.200 ;
        RECT 107.000 57.100 107.400 57.200 ;
        RECT 106.200 56.800 107.400 57.100 ;
        RECT 107.000 56.200 107.300 56.800 ;
        RECT 97.400 55.800 98.500 56.100 ;
        RECT 104.600 56.100 105.000 56.200 ;
        RECT 105.400 56.100 105.800 56.200 ;
        RECT 104.600 55.800 105.800 56.100 ;
        RECT 107.000 55.800 107.400 56.200 ;
        RECT 98.200 55.200 98.500 55.800 ;
        RECT 92.600 54.800 93.000 55.200 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 95.800 54.800 96.200 55.200 ;
        RECT 96.600 54.800 97.000 55.200 ;
        RECT 98.200 54.800 98.600 55.200 ;
        RECT 99.000 54.800 99.400 55.200 ;
        RECT 101.400 54.800 101.800 55.200 ;
        RECT 96.600 53.200 96.900 54.800 ;
        RECT 99.000 54.200 99.300 54.800 ;
        RECT 101.400 54.200 101.700 54.800 ;
        RECT 97.400 53.800 97.800 54.200 ;
        RECT 99.000 53.800 99.400 54.200 ;
        RECT 101.400 53.800 101.800 54.200 ;
        RECT 102.200 54.100 102.600 54.200 ;
        RECT 103.000 54.100 103.400 54.200 ;
        RECT 102.200 53.800 103.400 54.100 ;
        RECT 87.000 52.800 87.400 53.200 ;
        RECT 87.800 53.100 88.200 53.200 ;
        RECT 88.600 53.100 89.000 53.200 ;
        RECT 87.800 52.800 89.000 53.100 ;
        RECT 91.800 52.800 92.200 53.200 ;
        RECT 96.600 52.800 97.000 53.200 ;
        RECT 87.000 52.200 87.300 52.800 ;
        RECT 87.000 51.800 87.400 52.200 ;
        RECT 89.400 52.100 89.800 52.200 ;
        RECT 90.200 52.100 90.600 52.200 ;
        RECT 89.400 51.800 90.600 52.100 ;
        RECT 96.600 51.800 97.000 52.200 ;
        RECT 96.600 51.200 96.900 51.800 ;
        RECT 87.000 50.800 87.400 51.200 ;
        RECT 92.600 50.800 93.000 51.200 ;
        RECT 96.600 50.800 97.000 51.200 ;
        RECT 87.000 49.200 87.300 50.800 ;
        RECT 92.600 49.200 92.900 50.800 ;
        RECT 87.000 48.800 87.400 49.200 ;
        RECT 92.600 48.800 93.000 49.200 ;
        RECT 86.200 48.100 86.600 48.200 ;
        RECT 87.000 48.100 87.400 48.200 ;
        RECT 88.600 48.100 89.000 48.200 ;
        RECT 86.200 47.800 89.000 48.100 ;
        RECT 94.200 47.800 94.600 48.200 ;
        RECT 94.200 47.200 94.500 47.800 ;
        RECT 97.400 47.200 97.700 53.800 ;
        RECT 100.600 53.100 101.000 53.200 ;
        RECT 101.400 53.100 101.800 53.200 ;
        RECT 100.600 52.800 101.800 53.100 ;
        RECT 103.800 52.800 104.200 53.200 ;
        RECT 99.800 52.100 100.200 52.200 ;
        RECT 99.000 51.800 100.200 52.100 ;
        RECT 98.200 49.800 98.600 50.200 ;
        RECT 98.200 49.200 98.500 49.800 ;
        RECT 98.200 48.800 98.600 49.200 ;
        RECT 98.200 47.200 98.500 48.800 ;
        RECT 99.000 48.200 99.300 51.800 ;
        RECT 103.800 49.200 104.100 52.800 ;
        RECT 105.400 52.200 105.700 55.800 ;
        RECT 107.800 55.200 108.100 57.800 ;
        RECT 108.600 56.200 108.900 58.800 ;
        RECT 108.600 55.800 109.000 56.200 ;
        RECT 109.400 55.200 109.700 58.800 ;
        RECT 110.200 57.800 110.600 58.200 ;
        RECT 107.800 54.800 108.200 55.200 ;
        RECT 109.400 54.800 109.800 55.200 ;
        RECT 110.200 54.200 110.500 57.800 ;
        RECT 111.800 56.800 112.200 57.200 ;
        RECT 107.800 53.800 108.200 54.200 ;
        RECT 110.200 53.800 110.600 54.200 ;
        RECT 107.800 53.200 108.100 53.800 ;
        RECT 111.800 53.200 112.100 56.800 ;
        RECT 112.600 56.200 112.900 58.800 ;
        RECT 115.000 58.200 115.300 61.800 ;
        RECT 113.400 57.800 113.800 58.200 ;
        RECT 115.000 57.800 115.400 58.200 ;
        RECT 112.600 55.800 113.000 56.200 ;
        RECT 113.400 55.200 113.700 57.800 ;
        RECT 114.200 57.100 114.600 57.200 ;
        RECT 115.000 57.100 115.400 57.200 ;
        RECT 114.200 56.800 115.400 57.100 ;
        RECT 116.600 56.800 117.000 57.200 ;
        RECT 113.400 54.800 113.800 55.200 ;
        RECT 114.200 54.800 114.600 55.200 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 111.800 52.800 112.200 53.200 ;
        RECT 105.400 51.800 105.800 52.200 ;
        RECT 111.000 51.800 111.400 52.200 ;
        RECT 111.000 51.200 111.300 51.800 ;
        RECT 111.000 50.800 111.400 51.200 ;
        RECT 111.800 49.800 112.200 50.200 ;
        RECT 103.000 48.800 103.400 49.200 ;
        RECT 103.800 48.800 104.200 49.200 ;
        RECT 107.800 48.800 108.200 49.200 ;
        RECT 103.000 48.200 103.300 48.800 ;
        RECT 99.000 47.800 99.400 48.200 ;
        RECT 100.600 47.800 101.000 48.200 ;
        RECT 103.000 47.800 103.400 48.200 ;
        RECT 107.000 47.800 107.400 48.200 ;
        RECT 100.600 47.200 100.900 47.800 ;
        RECT 107.000 47.200 107.300 47.800 ;
        RECT 107.800 47.200 108.100 48.800 ;
        RECT 111.000 47.800 111.400 48.200 ;
        RECT 111.000 47.200 111.300 47.800 ;
        RECT 86.200 46.800 86.600 47.200 ;
        RECT 90.200 46.800 90.600 47.200 ;
        RECT 94.200 46.800 94.600 47.200 ;
        RECT 97.400 46.800 97.800 47.200 ;
        RECT 98.200 46.800 98.600 47.200 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 107.000 46.800 107.400 47.200 ;
        RECT 107.800 46.800 108.200 47.200 ;
        RECT 111.000 46.800 111.400 47.200 ;
        RECT 86.200 46.200 86.500 46.800 ;
        RECT 90.200 46.200 90.500 46.800 ;
        RECT 97.400 46.200 97.700 46.800 ;
        RECT 107.000 46.200 107.300 46.800 ;
        RECT 111.800 46.200 112.100 49.800 ;
        RECT 114.200 48.200 114.500 54.800 ;
        RECT 115.000 51.800 115.400 52.200 ;
        RECT 115.000 49.200 115.300 51.800 ;
        RECT 116.600 49.200 116.900 56.800 ;
        RECT 117.400 55.200 117.700 61.800 ;
        RECT 131.000 59.200 131.300 61.800 ;
        RECT 132.600 60.200 132.900 73.800 ;
        RECT 133.300 73.500 133.600 75.900 ;
        RECT 134.600 74.200 135.000 74.300 ;
        RECT 136.700 74.200 137.000 75.900 ;
        RECT 138.200 76.200 138.500 76.800 ;
        RECT 138.200 75.800 138.600 76.200 ;
        RECT 139.000 75.200 139.300 76.800 ;
        RECT 140.600 76.100 141.000 76.200 ;
        RECT 141.400 76.100 141.800 76.200 ;
        RECT 140.600 75.800 141.800 76.100 ;
        RECT 142.200 75.200 142.500 76.800 ;
        RECT 138.200 74.800 138.600 75.200 ;
        RECT 139.000 74.800 139.400 75.200 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 134.600 73.900 137.000 74.200 ;
        RECT 134.200 73.500 134.600 73.600 ;
        RECT 135.900 73.500 136.300 73.600 ;
        RECT 136.700 73.500 137.000 73.900 ;
        RECT 133.300 73.100 133.700 73.500 ;
        RECT 134.200 73.200 136.300 73.500 ;
        RECT 136.600 73.100 137.000 73.500 ;
        RECT 137.400 73.800 137.800 74.200 ;
        RECT 137.400 73.200 137.700 73.800 ;
        RECT 137.400 72.800 137.800 73.200 ;
        RECT 138.200 69.200 138.500 74.800 ;
        RECT 143.000 69.200 143.300 81.800 ;
        RECT 144.600 77.200 144.900 81.800 ;
        RECT 144.600 76.800 145.000 77.200 ;
        RECT 145.400 77.100 145.800 77.200 ;
        RECT 146.200 77.100 146.600 77.200 ;
        RECT 145.400 76.800 146.600 77.100 ;
        RECT 147.000 76.200 147.300 83.800 ;
        RECT 148.600 83.200 148.900 83.800 ;
        RECT 148.600 82.800 149.000 83.200 ;
        RECT 147.800 81.800 148.200 82.200 ;
        RECT 147.800 77.200 148.100 81.800 ;
        RECT 147.800 76.800 148.200 77.200 ;
        RECT 149.400 76.200 149.700 94.800 ;
        RECT 150.200 93.800 150.600 94.200 ;
        RECT 150.200 79.200 150.500 93.800 ;
        RECT 151.000 90.200 151.300 104.800 ;
        RECT 151.000 89.800 151.400 90.200 ;
        RECT 150.200 78.800 150.600 79.200 ;
        RECT 147.000 75.800 147.400 76.200 ;
        RECT 147.800 75.800 148.200 76.200 ;
        RECT 149.400 75.800 149.800 76.200 ;
        RECT 145.400 75.100 145.800 75.200 ;
        RECT 146.200 75.100 146.600 75.200 ;
        RECT 145.400 74.800 146.600 75.100 ;
        RECT 147.000 74.100 147.300 75.800 ;
        RECT 147.800 75.200 148.100 75.800 ;
        RECT 147.800 74.800 148.200 75.200 ;
        RECT 148.600 74.800 149.000 75.200 ;
        RECT 148.600 74.200 148.900 74.800 ;
        RECT 147.000 73.800 148.100 74.100 ;
        RECT 148.600 73.800 149.000 74.200 ;
        RECT 150.200 73.800 150.600 74.200 ;
        RECT 143.800 71.800 144.200 72.200 ;
        RECT 145.400 71.800 145.800 72.200 ;
        RECT 138.200 68.800 138.600 69.200 ;
        RECT 143.000 68.800 143.400 69.200 ;
        RECT 138.200 68.100 138.600 68.200 ;
        RECT 139.000 68.100 139.400 68.200 ;
        RECT 138.200 67.800 139.400 68.100 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 133.400 66.100 133.800 66.200 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 133.400 65.800 134.600 66.100 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 133.400 64.800 133.800 65.200 ;
        RECT 135.000 64.800 135.400 65.200 ;
        RECT 133.400 64.200 133.700 64.800 ;
        RECT 135.000 64.200 135.300 64.800 ;
        RECT 136.600 64.200 136.900 65.800 ;
        RECT 137.400 65.200 137.700 66.800 ;
        RECT 143.800 66.200 144.100 71.800 ;
        RECT 141.400 66.100 141.800 66.200 ;
        RECT 142.200 66.100 142.600 66.200 ;
        RECT 141.400 65.800 142.600 66.100 ;
        RECT 143.800 65.800 144.200 66.200 ;
        RECT 144.600 65.800 145.000 66.200 ;
        RECT 137.400 64.800 137.800 65.200 ;
        RECT 142.200 65.100 142.600 65.200 ;
        RECT 143.000 65.100 143.400 65.200 ;
        RECT 142.200 64.800 143.400 65.100 ;
        RECT 143.800 64.200 144.100 65.800 ;
        RECT 133.400 63.800 133.800 64.200 ;
        RECT 135.000 63.800 135.400 64.200 ;
        RECT 136.600 63.800 137.000 64.200 ;
        RECT 140.600 63.800 141.000 64.200 ;
        RECT 143.800 63.800 144.200 64.200 ;
        RECT 140.600 63.200 140.900 63.800 ;
        RECT 133.400 62.800 133.800 63.200 ;
        RECT 140.600 62.800 141.000 63.200 ;
        RECT 132.600 59.800 133.000 60.200 ;
        RECT 131.000 58.800 131.400 59.200 ;
        RECT 123.800 57.800 124.200 58.200 ;
        RECT 129.400 58.100 129.800 58.200 ;
        RECT 130.200 58.100 130.600 58.200 ;
        RECT 129.400 57.800 130.600 58.100 ;
        RECT 123.800 57.200 124.100 57.800 ;
        RECT 118.200 56.800 118.600 57.200 ;
        RECT 123.000 56.800 123.400 57.200 ;
        RECT 123.800 56.800 124.200 57.200 ;
        RECT 124.600 56.800 125.000 57.200 ;
        RECT 127.800 56.800 128.200 57.200 ;
        RECT 131.000 56.800 131.400 57.200 ;
        RECT 118.200 56.200 118.500 56.800 ;
        RECT 123.000 56.200 123.300 56.800 ;
        RECT 124.600 56.200 124.900 56.800 ;
        RECT 118.200 55.800 118.600 56.200 ;
        RECT 123.000 55.800 123.400 56.200 ;
        RECT 124.600 55.800 125.000 56.200 ;
        RECT 125.400 55.800 125.800 56.200 ;
        RECT 117.400 54.800 117.800 55.200 ;
        RECT 119.000 54.800 119.400 55.200 ;
        RECT 123.000 55.100 123.400 55.200 ;
        RECT 123.800 55.100 124.200 55.200 ;
        RECT 123.000 54.800 124.200 55.100 ;
        RECT 119.000 54.200 119.300 54.800 ;
        RECT 117.400 53.800 117.800 54.200 ;
        RECT 119.000 53.800 119.400 54.200 ;
        RECT 119.800 53.800 120.200 54.200 ;
        RECT 117.400 53.200 117.700 53.800 ;
        RECT 119.800 53.200 120.100 53.800 ;
        RECT 125.400 53.200 125.700 55.800 ;
        RECT 127.800 55.200 128.100 56.800 ;
        RECT 131.000 56.200 131.300 56.800 ;
        RECT 131.000 55.800 131.400 56.200 ;
        RECT 127.000 54.800 127.400 55.200 ;
        RECT 127.800 55.100 128.200 55.200 ;
        RECT 128.600 55.100 129.000 55.200 ;
        RECT 127.800 54.800 129.000 55.100 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 127.000 54.200 127.300 54.800 ;
        RECT 129.400 54.200 129.700 54.800 ;
        RECT 127.000 53.800 127.400 54.200 ;
        RECT 128.600 53.800 129.000 54.200 ;
        RECT 129.400 53.800 129.800 54.200 ;
        RECT 128.600 53.200 128.900 53.800 ;
        RECT 117.400 52.800 117.800 53.200 ;
        RECT 119.800 52.800 120.200 53.200 ;
        RECT 121.400 53.100 121.800 53.200 ;
        RECT 122.200 53.100 122.600 53.200 ;
        RECT 121.400 52.800 122.600 53.100 ;
        RECT 123.000 52.800 123.400 53.200 ;
        RECT 125.400 52.800 125.800 53.200 ;
        RECT 126.200 52.800 126.600 53.200 ;
        RECT 127.800 52.800 128.200 53.200 ;
        RECT 128.600 52.800 129.000 53.200 ;
        RECT 119.800 51.800 120.200 52.200 ;
        RECT 120.600 51.800 121.000 52.200 ;
        RECT 115.000 48.800 115.400 49.200 ;
        RECT 116.600 48.800 117.000 49.200 ;
        RECT 114.200 47.800 114.600 48.200 ;
        RECT 115.000 48.100 115.400 48.200 ;
        RECT 115.800 48.100 116.200 48.200 ;
        RECT 115.000 47.800 116.200 48.100 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 87.800 45.800 88.200 46.200 ;
        RECT 88.600 46.100 89.000 46.200 ;
        RECT 89.400 46.100 89.800 46.200 ;
        RECT 88.600 45.800 89.800 46.100 ;
        RECT 90.200 45.800 90.600 46.200 ;
        RECT 91.000 45.800 91.400 46.200 ;
        RECT 95.800 45.800 96.200 46.200 ;
        RECT 96.600 45.800 97.000 46.200 ;
        RECT 97.400 45.800 97.800 46.200 ;
        RECT 105.400 45.800 105.800 46.200 ;
        RECT 107.000 45.800 107.400 46.200 ;
        RECT 110.200 45.800 110.600 46.200 ;
        RECT 111.800 45.800 112.200 46.200 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 85.400 44.800 85.800 45.200 ;
        RECT 83.800 42.800 84.200 43.200 ;
        RECT 83.800 37.800 84.200 38.200 ;
        RECT 83.000 35.800 83.400 36.200 ;
        RECT 83.000 33.200 83.300 35.800 ;
        RECT 83.800 35.200 84.100 37.800 ;
        RECT 86.200 35.800 86.600 36.200 ;
        RECT 86.200 35.200 86.500 35.800 ;
        RECT 87.800 35.200 88.100 45.800 ;
        RECT 88.600 36.100 89.000 36.200 ;
        RECT 89.400 36.100 89.800 36.200 ;
        RECT 88.600 35.800 89.800 36.100 ;
        RECT 83.800 34.800 84.200 35.200 ;
        RECT 85.400 34.800 85.800 35.200 ;
        RECT 86.200 34.800 86.600 35.200 ;
        RECT 87.800 34.800 88.200 35.200 ;
        RECT 90.200 35.100 90.500 45.800 ;
        RECT 91.000 45.200 91.300 45.800 ;
        RECT 95.800 45.200 96.100 45.800 ;
        RECT 91.000 44.800 91.400 45.200 ;
        RECT 93.400 44.800 93.800 45.200 ;
        RECT 95.800 44.800 96.200 45.200 ;
        RECT 92.600 41.800 93.000 42.200 ;
        RECT 91.000 35.800 91.400 36.200 ;
        RECT 91.000 35.200 91.300 35.800 ;
        RECT 92.600 35.200 92.900 41.800 ;
        RECT 93.400 35.200 93.700 44.800 ;
        RECT 91.000 35.100 91.400 35.200 ;
        RECT 90.200 34.800 91.400 35.100 ;
        RECT 91.800 34.800 92.200 35.200 ;
        RECT 92.600 34.800 93.000 35.200 ;
        RECT 93.400 34.800 93.800 35.200 ;
        RECT 85.400 33.200 85.700 34.800 ;
        RECT 87.800 34.200 88.100 34.800 ;
        RECT 91.800 34.200 92.100 34.800 ;
        RECT 87.800 33.800 88.200 34.200 ;
        RECT 88.600 34.100 89.000 34.200 ;
        RECT 89.400 34.100 89.800 34.200 ;
        RECT 88.600 33.800 89.800 34.100 ;
        RECT 91.800 33.800 92.200 34.200 ;
        RECT 93.400 33.800 93.800 34.200 ;
        RECT 83.000 32.800 83.400 33.200 ;
        RECT 85.400 32.800 85.800 33.200 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 83.000 31.800 83.400 32.200 ;
        RECT 84.600 31.800 85.000 32.200 ;
        RECT 86.200 31.800 86.600 32.200 ;
        RECT 83.000 27.200 83.300 31.800 ;
        RECT 84.600 28.200 84.900 31.800 ;
        RECT 86.200 30.200 86.500 31.800 ;
        RECT 86.200 29.800 86.600 30.200 ;
        RECT 83.800 27.800 84.200 28.200 ;
        RECT 84.600 27.800 85.000 28.200 ;
        RECT 85.400 27.800 85.800 28.200 ;
        RECT 87.000 28.100 87.300 32.800 ;
        RECT 86.200 27.800 87.300 28.100 ;
        RECT 83.000 26.800 83.400 27.200 ;
        RECT 83.800 26.200 84.100 27.800 ;
        RECT 85.400 27.200 85.700 27.800 ;
        RECT 86.200 27.200 86.500 27.800 ;
        RECT 85.400 26.800 85.800 27.200 ;
        RECT 86.200 26.800 86.600 27.200 ;
        RECT 87.000 26.800 87.400 27.200 ;
        RECT 87.000 26.200 87.300 26.800 ;
        RECT 87.800 26.200 88.100 33.800 ;
        RECT 93.400 33.200 93.700 33.800 ;
        RECT 89.400 32.800 89.800 33.200 ;
        RECT 91.000 32.800 91.400 33.200 ;
        RECT 93.400 32.800 93.800 33.200 ;
        RECT 89.400 32.200 89.700 32.800 ;
        RECT 89.400 31.800 89.800 32.200 ;
        RECT 91.000 29.200 91.300 32.800 ;
        RECT 93.400 31.800 93.800 32.200 ;
        RECT 95.800 31.800 96.200 32.200 ;
        RECT 90.200 28.800 90.600 29.200 ;
        RECT 91.000 28.800 91.400 29.200 ;
        RECT 90.200 28.200 90.500 28.800 ;
        RECT 90.200 27.800 90.600 28.200 ;
        RECT 93.400 26.200 93.700 31.800 ;
        RECT 95.800 31.200 96.100 31.800 ;
        RECT 95.800 30.800 96.200 31.200 ;
        RECT 94.200 28.100 94.600 28.200 ;
        RECT 95.000 28.100 95.400 28.200 ;
        RECT 94.200 27.800 95.400 28.100 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 95.000 26.800 96.200 27.100 ;
        RECT 83.800 25.800 84.200 26.200 ;
        RECT 87.000 25.800 87.400 26.200 ;
        RECT 87.800 25.800 88.200 26.200 ;
        RECT 92.600 25.800 93.000 26.200 ;
        RECT 93.400 25.800 93.800 26.200 ;
        RECT 96.600 26.100 96.900 45.800 ;
        RECT 105.400 45.200 105.700 45.800 ;
        RECT 110.200 45.200 110.500 45.800 ;
        RECT 103.800 44.800 104.200 45.200 ;
        RECT 105.400 44.800 105.800 45.200 ;
        RECT 110.200 44.800 110.600 45.200 ;
        RECT 99.800 41.800 100.200 42.200 ;
        RECT 99.800 36.200 100.100 41.800 ;
        RECT 97.400 35.800 97.800 36.200 ;
        RECT 98.200 35.800 98.600 36.200 ;
        RECT 99.800 35.800 100.200 36.200 ;
        RECT 97.400 35.200 97.700 35.800 ;
        RECT 97.400 34.800 97.800 35.200 ;
        RECT 97.400 33.800 97.800 34.200 ;
        RECT 97.400 33.200 97.700 33.800 ;
        RECT 97.400 32.800 97.800 33.200 ;
        RECT 97.400 27.100 97.800 27.200 ;
        RECT 98.200 27.100 98.500 35.800 ;
        RECT 103.800 34.200 104.100 44.800 ;
        RECT 108.600 41.800 109.000 42.200 ;
        RECT 108.600 36.100 108.900 41.800 ;
        RECT 111.000 36.800 111.400 37.200 ;
        RECT 109.400 36.100 109.800 36.200 ;
        RECT 108.600 35.800 109.800 36.100 ;
        RECT 108.600 35.200 108.900 35.800 ;
        RECT 104.600 35.100 105.000 35.200 ;
        RECT 105.400 35.100 105.800 35.200 ;
        RECT 104.600 34.800 105.800 35.100 ;
        RECT 108.600 34.800 109.000 35.200 ;
        RECT 109.400 35.100 109.800 35.200 ;
        RECT 110.200 35.100 110.600 35.200 ;
        RECT 109.400 34.800 110.600 35.100 ;
        RECT 111.000 34.200 111.300 36.800 ;
        RECT 112.600 36.200 112.900 45.800 ;
        RECT 114.200 45.200 114.500 47.800 ;
        RECT 115.000 46.800 115.400 47.200 ;
        RECT 116.600 47.100 117.000 47.200 ;
        RECT 117.400 47.100 117.800 47.200 ;
        RECT 116.600 46.800 117.800 47.100 ;
        RECT 115.000 46.200 115.300 46.800 ;
        RECT 119.800 46.200 120.100 51.800 ;
        RECT 120.600 48.100 120.900 51.800 ;
        RECT 123.000 49.200 123.300 52.800 ;
        RECT 126.200 52.200 126.500 52.800 ;
        RECT 126.200 51.800 126.600 52.200 ;
        RECT 127.000 50.800 127.400 51.200 ;
        RECT 123.000 48.800 123.400 49.200 ;
        RECT 123.800 48.800 124.200 49.200 ;
        RECT 120.600 47.800 121.700 48.100 ;
        RECT 120.600 46.800 121.000 47.200 ;
        RECT 115.000 45.800 115.400 46.200 ;
        RECT 117.400 46.100 117.800 46.200 ;
        RECT 118.200 46.100 118.600 46.200 ;
        RECT 117.400 45.800 118.600 46.100 ;
        RECT 119.000 45.800 119.400 46.200 ;
        RECT 119.800 45.800 120.200 46.200 ;
        RECT 119.000 45.200 119.300 45.800 ;
        RECT 114.200 44.800 114.600 45.200 ;
        RECT 119.000 44.800 119.400 45.200 ;
        RECT 120.600 44.200 120.900 46.800 ;
        RECT 120.600 43.800 121.000 44.200 ;
        RECT 119.800 41.800 120.200 42.200 ;
        RECT 113.400 36.800 113.800 37.200 ;
        RECT 112.600 35.800 113.000 36.200 ;
        RECT 113.400 35.200 113.700 36.800 ;
        RECT 115.000 35.800 115.400 36.200 ;
        RECT 118.200 36.100 118.600 36.200 ;
        RECT 119.000 36.100 119.400 36.200 ;
        RECT 118.200 35.800 119.400 36.100 ;
        RECT 115.000 35.200 115.300 35.800 ;
        RECT 111.800 35.100 112.200 35.200 ;
        RECT 112.600 35.100 113.000 35.200 ;
        RECT 111.800 34.800 113.000 35.100 ;
        RECT 113.400 34.800 113.800 35.200 ;
        RECT 115.000 34.800 115.400 35.200 ;
        RECT 102.200 34.100 102.600 34.200 ;
        RECT 103.000 34.100 103.400 34.200 ;
        RECT 102.200 33.800 103.400 34.100 ;
        RECT 103.800 33.800 104.200 34.200 ;
        RECT 107.000 34.100 107.400 34.200 ;
        RECT 107.800 34.100 108.200 34.200 ;
        RECT 107.000 33.800 108.200 34.100 ;
        RECT 111.000 33.800 111.400 34.200 ;
        RECT 104.600 32.800 105.000 33.200 ;
        RECT 107.000 32.800 107.400 33.200 ;
        RECT 103.000 29.100 103.400 29.200 ;
        RECT 103.800 29.100 104.200 29.200 ;
        RECT 103.000 28.800 104.200 29.100 ;
        RECT 104.600 28.200 104.900 32.800 ;
        RECT 107.000 32.200 107.300 32.800 ;
        RECT 107.000 31.800 107.400 32.200 ;
        RECT 110.200 30.800 110.600 31.200 ;
        RECT 110.200 28.200 110.500 30.800 ;
        RECT 111.000 28.800 111.400 29.200 ;
        RECT 111.000 28.200 111.300 28.800 ;
        RECT 97.400 26.800 98.500 27.100 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 96.600 25.800 97.800 26.100 ;
        RECT 91.000 25.100 91.400 25.200 ;
        RECT 91.800 25.100 92.200 25.200 ;
        RECT 91.000 24.800 92.200 25.100 ;
        RECT 82.200 18.800 82.600 19.200 ;
        RECT 92.600 17.200 92.900 25.800 ;
        RECT 98.200 24.100 98.500 26.800 ;
        RECT 100.600 27.800 101.000 28.200 ;
        RECT 103.000 27.800 103.400 28.200 ;
        RECT 104.600 27.800 105.000 28.200 ;
        RECT 110.200 27.800 110.600 28.200 ;
        RECT 111.000 27.800 111.400 28.200 ;
        RECT 99.000 26.100 99.400 26.200 ;
        RECT 99.800 26.100 100.200 26.200 ;
        RECT 99.000 25.800 100.200 26.100 ;
        RECT 100.600 25.200 100.900 27.800 ;
        RECT 103.000 27.200 103.300 27.800 ;
        RECT 111.800 27.200 112.100 34.800 ;
        RECT 112.600 33.800 113.000 34.200 ;
        RECT 112.600 33.200 112.900 33.800 ;
        RECT 112.600 32.800 113.000 33.200 ;
        RECT 113.400 31.200 113.700 34.800 ;
        RECT 118.200 34.200 118.500 35.800 ;
        RECT 119.000 35.100 119.400 35.200 ;
        RECT 119.800 35.100 120.100 41.800 ;
        RECT 119.000 34.800 120.100 35.100 ;
        RECT 118.200 33.800 118.600 34.200 ;
        RECT 119.800 34.100 120.100 34.800 ;
        RECT 121.400 34.200 121.700 47.800 ;
        RECT 122.200 46.800 122.600 47.200 ;
        RECT 122.200 44.200 122.500 46.800 ;
        RECT 123.800 46.200 124.100 48.800 ;
        RECT 126.200 47.800 126.600 48.200 ;
        RECT 124.600 47.100 125.000 47.200 ;
        RECT 125.400 47.100 125.800 47.200 ;
        RECT 124.600 46.800 125.800 47.100 ;
        RECT 123.800 45.800 124.200 46.200 ;
        RECT 126.200 44.200 126.500 47.800 ;
        RECT 127.000 47.200 127.300 50.800 ;
        RECT 127.000 46.800 127.400 47.200 ;
        RECT 127.800 46.200 128.100 52.800 ;
        RECT 127.800 45.800 128.200 46.200 ;
        RECT 128.600 45.800 129.000 46.200 ;
        RECT 122.200 43.800 122.600 44.200 ;
        RECT 126.200 43.800 126.600 44.200 ;
        RECT 126.200 41.800 126.600 42.200 ;
        RECT 123.800 36.100 124.200 36.200 ;
        RECT 124.600 36.100 125.000 36.200 ;
        RECT 123.800 35.800 125.000 36.100 ;
        RECT 126.200 35.200 126.500 41.800 ;
        RECT 128.600 37.200 128.900 45.800 ;
        RECT 129.400 45.200 129.700 53.800 ;
        RECT 131.000 47.200 131.300 55.800 ;
        RECT 133.400 55.200 133.700 62.800 ;
        RECT 134.200 61.800 134.600 62.200 ;
        RECT 139.800 61.800 140.200 62.200 ;
        RECT 143.000 61.800 143.400 62.200 ;
        RECT 134.200 55.200 134.500 61.800 ;
        RECT 139.800 61.100 140.100 61.800 ;
        RECT 139.000 60.800 140.100 61.100 ;
        RECT 135.800 57.800 136.200 58.200 ;
        RECT 135.000 56.800 135.400 57.200 ;
        RECT 135.000 56.200 135.300 56.800 ;
        RECT 135.000 55.800 135.400 56.200 ;
        RECT 135.800 55.200 136.100 57.800 ;
        RECT 136.600 57.100 137.000 57.200 ;
        RECT 137.400 57.100 137.800 57.200 ;
        RECT 136.600 56.800 137.800 57.100 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 134.200 54.800 134.600 55.200 ;
        RECT 135.800 54.800 136.200 55.200 ;
        RECT 133.400 54.100 133.700 54.800 ;
        RECT 133.400 53.800 134.500 54.100 ;
        RECT 131.800 52.100 132.200 52.200 ;
        RECT 132.600 52.100 133.000 52.200 ;
        RECT 131.800 51.800 133.000 52.100 ;
        RECT 133.400 50.800 133.800 51.200 ;
        RECT 131.800 48.800 132.200 49.200 ;
        RECT 131.000 46.800 131.400 47.200 ;
        RECT 129.400 44.800 129.800 45.200 ;
        RECT 131.000 44.200 131.300 46.800 ;
        RECT 131.800 46.200 132.100 48.800 ;
        RECT 133.400 48.200 133.700 50.800 ;
        RECT 134.200 49.200 134.500 53.800 ;
        RECT 138.200 53.800 138.600 54.200 ;
        RECT 138.200 53.200 138.500 53.800 ;
        RECT 138.200 52.800 138.600 53.200 ;
        RECT 137.400 51.800 137.800 52.200 ;
        RECT 137.400 49.200 137.700 51.800 ;
        RECT 134.200 48.800 134.600 49.200 ;
        RECT 135.000 48.800 135.400 49.200 ;
        RECT 137.400 48.800 137.800 49.200 ;
        RECT 133.400 47.800 133.800 48.200 ;
        RECT 135.000 47.200 135.300 48.800 ;
        RECT 136.600 47.800 137.000 48.200 ;
        RECT 135.000 46.800 135.400 47.200 ;
        RECT 136.600 46.200 136.900 47.800 ;
        RECT 137.400 47.100 137.800 47.200 ;
        RECT 138.200 47.100 138.600 47.200 ;
        RECT 137.400 46.800 138.600 47.100 ;
        RECT 131.800 45.800 132.200 46.200 ;
        RECT 135.800 45.800 136.200 46.200 ;
        RECT 136.600 45.800 137.000 46.200 ;
        RECT 137.400 45.800 137.800 46.200 ;
        RECT 132.600 44.800 133.000 45.200 ;
        RECT 132.600 44.200 132.900 44.800 ;
        RECT 135.800 44.200 136.100 45.800 ;
        RECT 131.000 43.800 131.400 44.200 ;
        RECT 132.600 43.800 133.000 44.200 ;
        RECT 135.800 43.800 136.200 44.200 ;
        RECT 130.200 41.800 130.600 42.200 ;
        RECT 131.800 41.800 132.200 42.200 ;
        RECT 135.800 41.800 136.200 42.200 ;
        RECT 128.600 36.800 129.000 37.200 ;
        RECT 130.200 36.200 130.500 41.800 ;
        RECT 130.200 35.800 130.600 36.200 ;
        RECT 131.000 35.800 131.400 36.200 ;
        RECT 122.200 35.100 122.600 35.200 ;
        RECT 123.000 35.100 123.400 35.200 ;
        RECT 122.200 34.800 123.400 35.100 ;
        RECT 126.200 34.800 126.600 35.200 ;
        RECT 127.800 34.800 128.200 35.200 ;
        RECT 128.600 34.800 129.000 35.200 ;
        RECT 120.600 34.100 121.000 34.200 ;
        RECT 119.800 33.800 121.000 34.100 ;
        RECT 121.400 33.800 121.800 34.200 ;
        RECT 116.600 31.800 117.000 32.200 ;
        RECT 119.000 31.800 119.400 32.200 ;
        RECT 113.400 30.800 113.800 31.200 ;
        RECT 114.200 29.800 114.600 30.200 ;
        RECT 112.600 28.100 113.000 28.200 ;
        RECT 113.400 28.100 113.800 28.200 ;
        RECT 112.600 27.800 113.800 28.100 ;
        RECT 103.000 26.800 103.400 27.200 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 107.800 26.800 108.200 27.200 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 104.600 25.200 104.900 26.800 ;
        RECT 107.800 26.200 108.100 26.800 ;
        RECT 112.600 26.200 112.900 27.800 ;
        RECT 114.200 27.200 114.500 29.800 ;
        RECT 116.600 29.200 116.900 31.800 ;
        RECT 115.000 28.800 115.400 29.200 ;
        RECT 116.600 28.800 117.000 29.200 ;
        RECT 114.200 26.800 114.600 27.200 ;
        RECT 105.400 26.100 105.800 26.200 ;
        RECT 106.200 26.100 106.600 26.200 ;
        RECT 105.400 25.800 106.600 26.100 ;
        RECT 107.800 25.800 108.200 26.200 ;
        RECT 108.600 26.100 109.000 26.200 ;
        RECT 109.400 26.100 109.800 26.200 ;
        RECT 108.600 25.800 109.800 26.100 ;
        RECT 110.200 25.800 110.600 26.200 ;
        RECT 112.600 25.800 113.000 26.200 ;
        RECT 99.800 24.800 100.200 25.200 ;
        RECT 100.600 24.800 101.000 25.200 ;
        RECT 104.600 24.800 105.000 25.200 ;
        RECT 107.000 24.800 107.400 25.200 ;
        RECT 99.000 24.100 99.400 24.200 ;
        RECT 98.200 23.800 99.400 24.100 ;
        RECT 99.800 23.200 100.100 24.800 ;
        RECT 107.000 24.200 107.300 24.800 ;
        RECT 107.000 23.800 107.400 24.200 ;
        RECT 99.800 22.800 100.200 23.200 ;
        RECT 106.200 21.800 106.600 22.200 ;
        RECT 105.400 19.800 105.800 20.200 ;
        RECT 104.600 18.800 105.000 19.200 ;
        RECT 104.600 18.200 104.900 18.800 ;
        RECT 104.600 17.800 105.000 18.200 ;
        RECT 92.600 16.800 93.000 17.200 ;
        RECT 95.000 17.100 95.400 17.200 ;
        RECT 95.800 17.100 96.200 17.200 ;
        RECT 95.000 16.800 96.200 17.100 ;
        RECT 102.200 16.800 102.600 17.200 ;
        RECT 103.000 17.100 103.400 17.200 ;
        RECT 103.800 17.100 104.200 17.200 ;
        RECT 103.000 16.800 104.200 17.100 ;
        RECT 76.600 15.800 77.000 16.200 ;
        RECT 79.800 15.800 80.200 16.200 ;
        RECT 85.400 15.800 85.800 16.200 ;
        RECT 77.400 15.100 77.800 15.200 ;
        RECT 78.200 15.100 78.600 15.200 ;
        RECT 77.400 14.800 78.600 15.100 ;
        RECT 82.200 14.800 82.600 15.200 ;
        RECT 83.800 15.100 84.200 15.200 ;
        RECT 84.600 15.100 85.000 15.200 ;
        RECT 83.800 14.800 85.000 15.100 ;
        RECT 82.200 14.200 82.500 14.800 ;
        RECT 85.400 14.200 85.700 15.800 ;
        RECT 76.600 14.100 77.000 14.200 ;
        RECT 77.400 14.100 77.800 14.200 ;
        RECT 76.600 13.800 77.800 14.100 ;
        RECT 82.200 13.800 82.600 14.200 ;
        RECT 85.400 13.800 85.800 14.200 ;
        RECT 87.800 14.000 88.200 14.400 ;
        RECT 92.600 14.200 92.900 16.800 ;
        RECT 102.200 16.200 102.500 16.800 ;
        RECT 105.400 16.200 105.700 19.800 ;
        RECT 106.200 16.200 106.500 21.800 ;
        RECT 109.400 17.800 109.800 18.200 ;
        RECT 109.400 17.200 109.700 17.800 ;
        RECT 109.400 16.800 109.800 17.200 ;
        RECT 93.400 15.800 93.800 16.200 ;
        RECT 94.200 15.800 94.600 16.200 ;
        RECT 95.000 15.800 95.400 16.200 ;
        RECT 102.200 15.800 102.600 16.200 ;
        RECT 105.400 15.800 105.800 16.200 ;
        RECT 106.200 15.800 106.600 16.200 ;
        RECT 107.000 15.800 107.400 16.200 ;
        RECT 107.800 15.800 108.200 16.200 ;
        RECT 109.400 15.800 109.800 16.200 ;
        RECT 93.400 15.200 93.700 15.800 ;
        RECT 94.200 15.200 94.500 15.800 ;
        RECT 95.000 15.200 95.300 15.800 ;
        RECT 93.400 14.800 93.800 15.200 ;
        RECT 94.200 14.800 94.600 15.200 ;
        RECT 95.000 14.800 95.400 15.200 ;
        RECT 97.400 14.800 97.800 15.200 ;
        RECT 104.600 15.100 105.000 15.200 ;
        RECT 105.400 15.100 105.800 15.200 ;
        RECT 106.200 15.100 106.600 15.200 ;
        RECT 104.600 14.800 106.600 15.100 ;
        RECT 97.400 14.200 97.700 14.800 ;
        RECT 85.400 13.200 85.700 13.800 ;
        RECT 79.800 12.800 80.200 13.200 ;
        RECT 82.200 13.100 82.600 13.200 ;
        RECT 83.000 13.100 83.400 13.200 ;
        RECT 82.200 12.800 83.400 13.100 ;
        RECT 85.400 12.800 85.800 13.200 ;
        RECT 79.800 12.200 80.100 12.800 ;
        RECT 87.800 12.200 88.100 14.000 ;
        RECT 90.200 13.800 90.600 14.200 ;
        RECT 91.800 13.800 92.200 14.200 ;
        RECT 92.600 13.800 93.000 14.200 ;
        RECT 97.400 13.800 97.800 14.200 ;
        RECT 102.200 13.800 102.600 14.200 ;
        RECT 90.200 13.200 90.500 13.800 ;
        RECT 91.800 13.200 92.100 13.800 ;
        RECT 102.200 13.200 102.500 13.800 ;
        RECT 107.000 13.200 107.300 15.800 ;
        RECT 107.800 14.200 108.100 15.800 ;
        RECT 109.400 15.200 109.700 15.800 ;
        RECT 110.200 15.200 110.500 25.800 ;
        RECT 111.000 18.800 111.400 19.200 ;
        RECT 109.400 14.800 109.800 15.200 ;
        RECT 110.200 14.800 110.600 15.200 ;
        RECT 110.200 14.200 110.500 14.800 ;
        RECT 111.000 14.200 111.300 18.800 ;
        RECT 111.800 16.800 112.200 17.200 ;
        RECT 111.800 15.200 112.100 16.800 ;
        RECT 115.000 16.200 115.300 28.800 ;
        RECT 119.000 28.200 119.300 31.800 ;
        RECT 121.400 28.200 121.700 33.800 ;
        RECT 119.000 27.800 119.400 28.200 ;
        RECT 121.400 27.800 121.800 28.200 ;
        RECT 116.600 27.100 117.000 27.200 ;
        RECT 117.400 27.100 117.800 27.200 ;
        RECT 116.600 26.800 117.800 27.100 ;
        RECT 119.000 26.800 119.400 27.200 ;
        RECT 119.800 27.100 120.200 27.200 ;
        RECT 120.600 27.100 121.000 27.200 ;
        RECT 119.800 26.800 121.000 27.100 ;
        RECT 119.000 24.200 119.300 26.800 ;
        RECT 123.000 26.200 123.300 34.800 ;
        RECT 123.800 34.100 124.200 34.200 ;
        RECT 124.600 34.100 125.000 34.200 ;
        RECT 123.800 33.800 125.000 34.100 ;
        RECT 125.400 34.100 125.800 34.200 ;
        RECT 126.200 34.100 126.600 34.200 ;
        RECT 125.400 33.800 126.600 34.100 ;
        RECT 124.600 32.800 125.000 33.200 ;
        RECT 125.400 32.800 125.800 33.200 ;
        RECT 123.000 25.800 123.400 26.200 ;
        RECT 119.000 23.800 119.400 24.200 ;
        RECT 115.800 21.800 116.200 22.200 ;
        RECT 115.800 20.200 116.100 21.800 ;
        RECT 115.800 19.800 116.200 20.200 ;
        RECT 124.600 19.200 124.900 32.800 ;
        RECT 125.400 32.200 125.700 32.800 ;
        RECT 125.400 31.800 125.800 32.200 ;
        RECT 125.400 28.100 125.800 28.200 ;
        RECT 126.200 28.100 126.600 28.200 ;
        RECT 125.400 27.800 126.600 28.100 ;
        RECT 127.000 27.800 127.400 28.200 ;
        RECT 125.400 26.800 125.800 27.200 ;
        RECT 125.400 25.200 125.700 26.800 ;
        RECT 126.200 25.800 126.600 26.200 ;
        RECT 125.400 24.800 125.800 25.200 ;
        RECT 124.600 18.800 125.000 19.200 ;
        RECT 126.200 17.200 126.500 25.800 ;
        RECT 122.200 16.800 122.600 17.200 ;
        RECT 126.200 16.800 126.600 17.200 ;
        RECT 115.000 15.800 115.400 16.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 115.000 14.200 115.300 15.800 ;
        RECT 115.800 15.100 116.200 15.200 ;
        RECT 116.600 15.100 117.000 15.200 ;
        RECT 115.800 14.800 117.000 15.100 ;
        RECT 122.200 14.200 122.500 16.800 ;
        RECT 125.400 15.800 125.800 16.200 ;
        RECT 126.200 15.800 126.600 16.200 ;
        RECT 125.400 15.200 125.700 15.800 ;
        RECT 123.000 15.100 123.400 15.200 ;
        RECT 123.800 15.100 124.200 15.200 ;
        RECT 123.000 14.800 124.200 15.100 ;
        RECT 125.400 14.800 125.800 15.200 ;
        RECT 126.200 14.200 126.500 15.800 ;
        RECT 127.000 15.200 127.300 27.800 ;
        RECT 127.800 26.200 128.100 34.800 ;
        RECT 128.600 27.200 128.900 34.800 ;
        RECT 131.000 29.200 131.300 35.800 ;
        RECT 131.800 35.200 132.100 41.800 ;
        RECT 133.400 35.800 133.800 36.200 ;
        RECT 133.400 35.200 133.700 35.800 ;
        RECT 131.800 34.800 132.200 35.200 ;
        RECT 133.400 34.800 133.800 35.200 ;
        RECT 129.400 28.800 129.800 29.200 ;
        RECT 131.000 28.800 131.400 29.200 ;
        RECT 129.400 27.200 129.700 28.800 ;
        RECT 133.400 28.200 133.700 34.800 ;
        RECT 135.800 34.200 136.100 41.800 ;
        RECT 136.600 35.800 137.000 36.200 ;
        RECT 136.600 35.200 136.900 35.800 ;
        RECT 136.600 34.800 137.000 35.200 ;
        RECT 134.200 33.800 134.600 34.200 ;
        RECT 135.800 33.800 136.200 34.200 ;
        RECT 134.200 33.200 134.500 33.800 ;
        RECT 134.200 32.800 134.600 33.200 ;
        RECT 134.200 28.200 134.500 32.800 ;
        RECT 133.400 27.800 133.800 28.200 ;
        RECT 134.200 27.800 134.600 28.200 ;
        RECT 128.600 26.800 129.000 27.200 ;
        RECT 129.400 26.800 129.800 27.200 ;
        RECT 131.000 27.100 131.400 27.200 ;
        RECT 131.800 27.100 132.200 27.200 ;
        RECT 131.000 26.800 132.200 27.100 ;
        RECT 136.600 26.800 137.000 27.200 ;
        RECT 129.400 26.200 129.700 26.800 ;
        RECT 136.600 26.200 136.900 26.800 ;
        RECT 127.800 25.800 128.200 26.200 ;
        RECT 129.400 25.800 129.800 26.200 ;
        RECT 131.000 25.800 131.400 26.200 ;
        RECT 131.800 25.800 132.200 26.200 ;
        RECT 132.600 26.100 133.000 26.200 ;
        RECT 133.400 26.100 133.800 26.200 ;
        RECT 132.600 25.800 133.800 26.100 ;
        RECT 134.200 25.800 134.600 26.200 ;
        RECT 136.600 25.800 137.000 26.200 ;
        RECT 131.000 25.200 131.300 25.800 ;
        RECT 131.800 25.200 132.100 25.800 ;
        RECT 131.000 24.800 131.400 25.200 ;
        RECT 131.800 24.800 132.200 25.200 ;
        RECT 128.600 21.800 129.000 22.200 ;
        RECT 128.600 19.200 128.900 21.800 ;
        RECT 128.600 18.800 129.000 19.200 ;
        RECT 132.600 16.800 133.000 17.200 ;
        RECT 130.200 15.900 130.600 16.300 ;
        RECT 127.000 14.800 127.400 15.200 ;
        RECT 130.200 14.200 130.500 15.900 ;
        RECT 132.600 15.200 132.900 16.800 ;
        RECT 133.500 15.900 133.900 16.300 ;
        RECT 132.600 14.800 133.000 15.200 ;
        RECT 132.200 14.200 132.600 14.300 ;
        RECT 107.800 13.800 108.200 14.200 ;
        RECT 110.200 13.800 110.600 14.200 ;
        RECT 111.000 13.800 111.400 14.200 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 115.000 13.800 115.400 14.200 ;
        RECT 120.600 13.800 121.000 14.200 ;
        RECT 122.200 13.800 122.600 14.200 ;
        RECT 126.200 13.800 126.600 14.200 ;
        RECT 130.200 13.900 132.600 14.200 ;
        RECT 114.200 13.200 114.500 13.800 ;
        RECT 120.600 13.200 120.900 13.800 ;
        RECT 130.200 13.500 130.500 13.900 ;
        RECT 130.900 13.500 131.300 13.600 ;
        RECT 132.600 13.500 133.000 13.600 ;
        RECT 133.600 13.500 133.900 15.900 ;
        RECT 134.200 14.200 134.500 25.800 ;
        RECT 137.400 25.200 137.700 45.800 ;
        RECT 138.200 41.800 138.600 42.200 ;
        RECT 138.200 37.200 138.500 41.800 ;
        RECT 138.200 36.800 138.600 37.200 ;
        RECT 139.000 36.200 139.300 60.800 ;
        RECT 139.800 59.800 140.200 60.200 ;
        RECT 139.800 56.200 140.100 59.800 ;
        RECT 143.000 59.200 143.300 61.800 ;
        RECT 143.000 58.800 143.400 59.200 ;
        RECT 144.600 58.200 144.900 65.800 ;
        RECT 145.400 65.200 145.700 71.800 ;
        RECT 147.800 69.200 148.100 73.800 ;
        RECT 150.200 73.200 150.500 73.800 ;
        RECT 150.200 72.800 150.600 73.200 ;
        RECT 147.800 68.800 148.200 69.200 ;
        RECT 146.200 67.800 146.600 68.200 ;
        RECT 146.200 67.200 146.500 67.800 ;
        RECT 147.000 67.500 147.400 67.900 ;
        RECT 150.100 67.800 150.500 67.900 ;
        RECT 147.700 67.500 150.500 67.800 ;
        RECT 146.200 66.800 146.600 67.200 ;
        RECT 147.000 67.100 147.300 67.500 ;
        RECT 147.700 67.400 148.100 67.500 ;
        RECT 149.400 67.400 149.800 67.500 ;
        RECT 147.000 66.800 149.800 67.100 ;
        RECT 145.400 64.800 145.800 65.200 ;
        RECT 147.000 65.100 147.300 66.800 ;
        RECT 149.500 66.100 149.800 66.800 ;
        RECT 149.500 65.700 149.900 66.100 ;
        RECT 150.200 65.100 150.500 67.500 ;
        RECT 147.000 64.700 147.400 65.100 ;
        RECT 150.100 64.700 150.500 65.100 ;
        RECT 151.000 66.800 151.400 67.200 ;
        RECT 149.400 61.800 149.800 62.200 ;
        RECT 147.000 58.800 147.400 59.200 ;
        RECT 144.600 57.800 145.000 58.200 ;
        RECT 139.800 55.800 140.200 56.200 ;
        RECT 143.000 55.900 143.400 56.300 ;
        RECT 146.300 55.900 146.700 56.300 ;
        RECT 139.800 54.800 140.200 55.200 ;
        RECT 139.800 54.200 140.100 54.800 ;
        RECT 143.000 54.200 143.300 55.900 ;
        RECT 145.000 54.200 145.400 54.300 ;
        RECT 139.800 53.800 140.200 54.200 ;
        RECT 140.600 54.100 141.000 54.200 ;
        RECT 141.400 54.100 141.800 54.200 ;
        RECT 140.600 53.800 141.800 54.100 ;
        RECT 143.000 53.900 145.400 54.200 ;
        RECT 143.000 53.500 143.300 53.900 ;
        RECT 143.700 53.500 144.100 53.600 ;
        RECT 145.400 53.500 145.800 53.600 ;
        RECT 146.400 53.500 146.700 55.900 ;
        RECT 143.000 53.100 143.400 53.500 ;
        RECT 143.700 53.200 145.800 53.500 ;
        RECT 146.300 53.100 146.700 53.500 ;
        RECT 147.000 54.200 147.300 58.800 ;
        RECT 148.600 57.800 149.000 58.200 ;
        RECT 148.600 57.200 148.900 57.800 ;
        RECT 148.600 56.800 149.000 57.200 ;
        RECT 149.400 56.100 149.700 61.800 ;
        RECT 151.000 60.200 151.300 66.800 ;
        RECT 151.000 59.800 151.400 60.200 ;
        RECT 150.200 56.100 150.600 56.200 ;
        RECT 149.400 55.800 150.600 56.100 ;
        RECT 147.800 55.100 148.200 55.200 ;
        RECT 148.600 55.100 149.000 55.200 ;
        RECT 147.800 54.800 149.000 55.100 ;
        RECT 149.400 54.800 149.800 55.200 ;
        RECT 147.000 53.800 147.400 54.200 ;
        RECT 147.800 54.100 148.200 54.200 ;
        RECT 148.600 54.100 149.000 54.200 ;
        RECT 147.800 53.800 149.000 54.100 ;
        RECT 140.600 51.800 141.000 52.200 ;
        RECT 145.400 51.800 145.800 52.200 ;
        RECT 139.800 47.100 140.200 47.200 ;
        RECT 140.600 47.100 140.900 51.800 ;
        RECT 145.400 49.200 145.700 51.800 ;
        RECT 145.400 48.800 145.800 49.200 ;
        RECT 139.800 46.800 140.900 47.100 ;
        RECT 145.400 47.800 145.800 48.200 ;
        RECT 145.400 47.200 145.700 47.800 ;
        RECT 147.000 47.200 147.300 53.800 ;
        RECT 145.400 46.800 145.800 47.200 ;
        RECT 147.000 46.800 147.400 47.200 ;
        RECT 148.600 46.800 149.000 47.200 ;
        RECT 147.000 46.200 147.300 46.800 ;
        RECT 148.600 46.200 148.900 46.800 ;
        RECT 139.800 45.800 140.200 46.200 ;
        RECT 141.400 45.800 141.800 46.200 ;
        RECT 143.000 45.800 143.400 46.200 ;
        RECT 147.000 45.800 147.400 46.200 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 139.800 45.200 140.100 45.800 ;
        RECT 141.400 45.200 141.700 45.800 ;
        RECT 143.000 45.200 143.300 45.800 ;
        RECT 139.800 44.800 140.200 45.200 ;
        RECT 141.400 44.800 141.800 45.200 ;
        RECT 143.000 44.800 143.400 45.200 ;
        RECT 143.800 44.100 144.200 44.200 ;
        RECT 144.600 44.100 145.000 44.200 ;
        RECT 143.800 43.800 145.000 44.100 ;
        RECT 147.000 43.800 147.400 44.200 ;
        RECT 147.800 43.800 148.200 44.200 ;
        RECT 143.000 41.800 143.400 42.200 ;
        RECT 139.000 35.800 139.400 36.200 ;
        RECT 143.000 36.100 143.300 41.800 ;
        RECT 145.400 37.100 145.800 37.200 ;
        RECT 146.200 37.100 146.600 37.200 ;
        RECT 145.400 36.800 146.600 37.100 ;
        RECT 147.000 36.200 147.300 43.800 ;
        RECT 143.800 36.100 144.200 36.200 ;
        RECT 143.000 35.800 144.200 36.100 ;
        RECT 147.000 35.800 147.400 36.200 ;
        RECT 138.200 35.100 138.600 35.200 ;
        RECT 139.000 35.100 139.400 35.200 ;
        RECT 138.200 34.800 139.400 35.100 ;
        RECT 140.600 34.800 141.000 35.200 ;
        RECT 143.000 34.800 143.400 35.200 ;
        RECT 143.800 35.100 144.200 35.200 ;
        RECT 144.600 35.100 145.000 35.200 ;
        RECT 143.800 34.800 145.000 35.100 ;
        RECT 147.800 35.100 148.100 43.800 ;
        RECT 148.600 35.100 149.000 35.200 ;
        RECT 147.800 34.800 149.000 35.100 ;
        RECT 140.600 34.200 140.900 34.800 ;
        RECT 143.000 34.200 143.300 34.800 ;
        RECT 139.000 33.800 139.400 34.200 ;
        RECT 140.600 33.800 141.000 34.200 ;
        RECT 141.400 33.800 141.800 34.200 ;
        RECT 143.000 33.800 143.400 34.200 ;
        RECT 139.000 33.200 139.300 33.800 ;
        RECT 139.000 32.800 139.400 33.200 ;
        RECT 141.400 32.200 141.700 33.800 ;
        RECT 142.200 33.100 142.600 33.200 ;
        RECT 143.000 33.100 143.400 33.200 ;
        RECT 142.200 32.800 143.400 33.100 ;
        RECT 141.400 31.800 141.800 32.200 ;
        RECT 145.400 31.800 145.800 32.200 ;
        RECT 147.000 31.800 147.400 32.200 ;
        RECT 144.600 30.800 145.000 31.200 ;
        RECT 138.200 26.800 138.600 27.200 ;
        RECT 143.000 27.100 143.400 27.200 ;
        RECT 143.800 27.100 144.200 27.200 ;
        RECT 143.000 26.800 144.200 27.100 ;
        RECT 138.200 26.200 138.500 26.800 ;
        RECT 144.600 26.200 144.900 30.800 ;
        RECT 145.400 27.200 145.700 31.800 ;
        RECT 147.000 31.200 147.300 31.800 ;
        RECT 147.000 30.800 147.400 31.200 ;
        RECT 147.000 29.800 147.400 30.200 ;
        RECT 147.000 29.200 147.300 29.800 ;
        RECT 147.000 28.800 147.400 29.200 ;
        RECT 145.400 26.800 145.800 27.200 ;
        RECT 138.200 25.800 138.600 26.200 ;
        RECT 139.000 25.800 139.400 26.200 ;
        RECT 139.800 25.800 140.200 26.200 ;
        RECT 144.600 25.800 145.000 26.200 ;
        RECT 137.400 24.800 137.800 25.200 ;
        RECT 135.000 24.100 135.400 24.200 ;
        RECT 135.800 24.100 136.200 24.200 ;
        RECT 135.000 23.800 136.200 24.100 ;
        RECT 136.600 23.800 137.000 24.200 ;
        RECT 136.600 23.200 136.900 23.800 ;
        RECT 136.600 22.800 137.000 23.200 ;
        RECT 139.000 22.200 139.300 25.800 ;
        RECT 139.800 25.200 140.100 25.800 ;
        RECT 139.800 24.800 140.200 25.200 ;
        RECT 140.600 24.800 141.000 25.200 ;
        RECT 141.400 24.800 141.800 25.200 ;
        RECT 143.000 25.100 143.400 25.200 ;
        RECT 143.800 25.100 144.200 25.200 ;
        RECT 143.000 24.800 144.200 25.100 ;
        RECT 146.200 25.100 146.600 25.200 ;
        RECT 147.000 25.100 147.400 25.200 ;
        RECT 146.200 24.800 147.400 25.100 ;
        RECT 140.600 23.200 140.900 24.800 ;
        RECT 141.400 24.200 141.700 24.800 ;
        RECT 141.400 23.800 141.800 24.200 ;
        RECT 144.600 23.800 145.000 24.200 ;
        RECT 145.400 23.800 145.800 24.200 ;
        RECT 144.600 23.200 144.900 23.800 ;
        RECT 140.600 22.800 141.000 23.200 ;
        RECT 144.600 22.800 145.000 23.200 ;
        RECT 139.000 21.800 139.400 22.200 ;
        RECT 142.200 21.800 142.600 22.200 ;
        RECT 134.200 13.800 134.600 14.200 ;
        RECT 90.200 12.800 90.600 13.200 ;
        RECT 91.800 12.800 92.200 13.200 ;
        RECT 96.600 13.100 97.000 13.200 ;
        RECT 97.400 13.100 97.800 13.200 ;
        RECT 96.600 12.800 97.800 13.100 ;
        RECT 102.200 12.800 102.600 13.200 ;
        RECT 107.000 12.800 107.400 13.200 ;
        RECT 114.200 12.800 114.600 13.200 ;
        RECT 120.600 12.800 121.000 13.200 ;
        RECT 121.400 12.800 121.800 13.200 ;
        RECT 123.000 13.100 123.400 13.200 ;
        RECT 123.800 13.100 124.200 13.200 ;
        RECT 130.200 13.100 130.600 13.500 ;
        RECT 130.900 13.200 133.000 13.500 ;
        RECT 133.500 13.100 133.900 13.500 ;
        RECT 135.000 13.100 135.400 15.900 ;
        RECT 135.800 13.800 136.200 14.200 ;
        RECT 123.000 12.800 124.200 13.100 ;
        RECT 121.400 12.200 121.700 12.800 ;
        RECT 79.800 11.800 80.200 12.200 ;
        RECT 83.000 11.800 83.400 12.200 ;
        RECT 86.200 11.800 86.600 12.200 ;
        RECT 87.800 11.800 88.200 12.200 ;
        RECT 98.200 11.800 98.600 12.200 ;
        RECT 113.400 11.800 113.800 12.200 ;
        RECT 121.400 11.800 121.800 12.200 ;
        RECT 124.600 11.800 125.000 12.200 ;
        RECT 83.000 10.100 83.300 11.800 ;
        RECT 82.200 9.800 83.300 10.100 ;
        RECT 75.800 6.800 76.200 7.200 ;
        RECT 78.200 3.100 78.600 8.900 ;
        RECT 79.800 7.100 80.200 7.200 ;
        RECT 80.600 7.100 81.000 7.200 ;
        RECT 79.800 6.800 81.000 7.100 ;
        RECT 82.200 6.300 82.500 9.800 ;
        RECT 82.200 5.900 82.600 6.300 ;
        RECT 83.000 3.100 83.400 8.900 ;
        RECT 84.600 5.100 85.000 7.900 ;
        RECT 85.400 5.100 85.800 7.900 ;
        RECT 86.200 6.200 86.500 11.800 ;
        RECT 86.200 5.800 86.600 6.200 ;
        RECT 87.000 3.100 87.400 8.900 ;
        RECT 91.000 7.800 91.400 8.200 ;
        RECT 91.000 7.200 91.300 7.800 ;
        RECT 87.800 6.800 88.200 7.200 ;
        RECT 91.000 6.800 91.400 7.200 ;
        RECT 87.800 6.300 88.100 6.800 ;
        RECT 87.800 5.900 88.200 6.300 ;
        RECT 91.800 3.100 92.200 8.900 ;
        RECT 98.200 6.200 98.500 11.800 ;
        RECT 98.200 5.800 98.600 6.200 ;
        RECT 99.000 5.100 99.400 7.900 ;
        RECT 99.800 7.800 100.200 8.200 ;
        RECT 99.800 7.200 100.100 7.800 ;
        RECT 99.800 6.800 100.200 7.200 ;
        RECT 100.600 3.100 101.000 8.900 ;
        RECT 101.400 6.800 101.800 7.200 ;
        RECT 101.400 6.300 101.700 6.800 ;
        RECT 101.400 5.900 101.800 6.300 ;
        RECT 105.400 3.100 105.800 8.900 ;
        RECT 111.000 5.100 111.400 7.900 ;
        RECT 111.800 7.800 112.200 8.200 ;
        RECT 111.800 7.200 112.100 7.800 ;
        RECT 111.800 6.800 112.200 7.200 ;
        RECT 112.600 3.100 113.000 8.900 ;
        RECT 113.400 6.300 113.700 11.800 ;
        RECT 124.600 10.100 124.900 11.800 ;
        RECT 124.600 9.800 125.700 10.100 ;
        RECT 113.400 5.900 113.800 6.300 ;
        RECT 117.400 3.100 117.800 8.900 ;
        RECT 123.000 5.100 123.400 7.900 ;
        RECT 123.800 7.800 124.200 8.200 ;
        RECT 123.800 7.200 124.100 7.800 ;
        RECT 123.800 6.800 124.200 7.200 ;
        RECT 124.600 3.100 125.000 8.900 ;
        RECT 125.400 6.300 125.700 9.800 ;
        RECT 125.400 5.900 125.800 6.300 ;
        RECT 129.400 3.100 129.800 8.900 ;
        RECT 135.800 8.200 136.100 13.800 ;
        RECT 136.600 12.100 137.000 17.900 ;
        RECT 137.400 15.800 137.800 16.200 ;
        RECT 137.400 15.100 137.700 15.800 ;
        RECT 137.400 14.700 137.800 15.100 ;
        RECT 141.400 12.100 141.800 17.900 ;
        RECT 135.000 5.100 135.400 7.900 ;
        RECT 135.800 7.800 136.200 8.200 ;
        RECT 135.800 7.200 136.100 7.800 ;
        RECT 135.800 6.800 136.200 7.200 ;
        RECT 136.600 3.100 137.000 8.900 ;
        RECT 138.200 6.100 138.600 6.200 ;
        RECT 139.000 6.100 139.400 6.200 ;
        RECT 138.200 5.800 139.400 6.100 ;
        RECT 141.400 3.100 141.800 8.900 ;
        RECT 142.200 6.200 142.500 21.800 ;
        RECT 145.400 13.200 145.700 23.800 ;
        RECT 147.800 20.100 148.100 34.800 ;
        RECT 149.400 27.200 149.700 54.800 ;
        RECT 150.200 41.800 150.600 42.200 ;
        RECT 150.200 34.200 150.500 41.800 ;
        RECT 150.200 33.800 150.600 34.200 ;
        RECT 148.600 26.800 149.000 27.200 ;
        RECT 149.400 26.800 149.800 27.200 ;
        RECT 148.600 26.200 148.900 26.800 ;
        RECT 148.600 25.800 149.000 26.200 ;
        RECT 147.000 19.800 148.100 20.100 ;
        RECT 147.000 15.200 147.300 19.800 ;
        RECT 147.800 18.800 148.200 19.200 ;
        RECT 147.800 18.200 148.100 18.800 ;
        RECT 147.800 17.800 148.200 18.200 ;
        RECT 148.600 16.100 149.000 16.200 ;
        RECT 149.400 16.100 149.800 16.200 ;
        RECT 148.600 15.800 149.800 16.100 ;
        RECT 147.000 14.800 147.400 15.200 ;
        RECT 147.000 14.100 147.400 14.200 ;
        RECT 147.800 14.100 148.200 14.200 ;
        RECT 147.000 13.800 148.200 14.100 ;
        RECT 145.400 12.800 145.800 13.200 ;
        RECT 147.000 12.800 147.400 13.200 ;
        RECT 147.000 9.200 147.300 12.800 ;
        RECT 147.000 8.800 147.400 9.200 ;
        RECT 148.600 7.200 148.900 15.800 ;
        RECT 150.200 14.200 150.500 33.800 ;
        RECT 150.200 13.800 150.600 14.200 ;
        RECT 148.600 6.800 149.000 7.200 ;
        RECT 142.200 5.800 142.600 6.200 ;
        RECT 147.000 5.800 147.400 6.200 ;
        RECT 147.000 5.200 147.300 5.800 ;
        RECT 147.000 4.800 147.400 5.200 ;
      LAYER via2 ;
        RECT 30.200 128.800 30.600 129.200 ;
        RECT 1.400 127.800 1.800 128.200 ;
        RECT 11.000 126.800 11.400 127.200 ;
        RECT 14.200 125.800 14.600 126.200 ;
        RECT 20.600 126.800 21.000 127.200 ;
        RECT 17.400 115.800 17.800 116.200 ;
        RECT 20.600 108.800 21.000 109.200 ;
        RECT 15.800 87.800 16.200 88.200 ;
        RECT 19.000 85.800 19.400 86.200 ;
        RECT 2.200 71.800 2.600 72.200 ;
        RECT 39.800 114.800 40.200 115.200 ;
        RECT 39.800 112.800 40.200 113.200 ;
        RECT 39.000 111.800 39.400 112.200 ;
        RECT 36.600 106.800 37.000 107.200 ;
        RECT 36.600 104.800 37.000 105.200 ;
        RECT 59.800 114.800 60.200 115.200 ;
        RECT 55.000 113.800 55.400 114.200 ;
        RECT 48.600 106.800 49.000 107.200 ;
        RECT 39.000 94.800 39.400 95.200 ;
        RECT 37.400 92.800 37.800 93.200 ;
        RECT 31.800 65.800 32.200 66.200 ;
        RECT 31.800 58.800 32.200 59.200 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 48.600 85.800 49.000 86.200 ;
        RECT 48.600 71.800 49.000 72.200 ;
        RECT 65.400 101.800 65.800 102.200 ;
        RECT 63.800 93.800 64.200 94.200 ;
        RECT 63.800 92.800 64.200 93.200 ;
        RECT 59.000 81.800 59.400 82.200 ;
        RECT 92.600 125.800 93.000 126.200 ;
        RECT 87.800 115.800 88.200 116.200 ;
        RECT 72.600 111.800 73.000 112.200 ;
        RECT 71.000 94.800 71.400 95.200 ;
        RECT 70.200 93.800 70.600 94.200 ;
        RECT 81.400 106.800 81.800 107.200 ;
        RECT 98.200 113.800 98.600 114.200 ;
        RECT 89.400 104.800 89.800 105.200 ;
        RECT 88.600 102.800 89.000 103.200 ;
        RECT 85.400 98.800 85.800 99.200 ;
        RECT 122.200 125.800 122.600 126.200 ;
        RECT 147.800 127.800 148.200 128.200 ;
        RECT 125.400 123.800 125.800 124.200 ;
        RECT 128.600 123.800 129.000 124.200 ;
        RECT 135.000 122.800 135.400 123.200 ;
        RECT 79.800 96.800 80.200 97.200 ;
        RECT 93.400 96.800 93.800 97.200 ;
        RECT 83.800 94.800 84.200 95.200 ;
        RECT 60.600 76.800 61.000 77.200 ;
        RECT 62.200 75.800 62.600 76.200 ;
        RECT 83.000 86.800 83.400 87.200 ;
        RECT 89.400 95.800 89.800 96.200 ;
        RECT 96.600 95.800 97.000 96.200 ;
        RECT 75.000 74.800 75.400 75.200 ;
        RECT 59.000 55.800 59.400 56.200 ;
        RECT 62.200 53.800 62.600 54.200 ;
        RECT 101.400 93.800 101.800 94.200 ;
        RECT 98.200 86.800 98.600 87.200 ;
        RECT 96.600 81.800 97.000 82.200 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 75.000 53.800 75.400 54.200 ;
        RECT 79.800 65.800 80.200 66.200 ;
        RECT 80.600 63.800 81.000 64.200 ;
        RECT 35.000 47.800 35.400 48.200 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 35.000 45.800 35.400 46.200 ;
        RECT 38.200 45.800 38.600 46.200 ;
        RECT 14.200 11.800 14.600 12.200 ;
        RECT 43.000 44.800 43.400 45.200 ;
        RECT 67.800 45.800 68.200 46.200 ;
        RECT 51.800 28.800 52.200 29.200 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 63.000 28.800 63.400 29.200 ;
        RECT 7.000 6.800 7.400 7.200 ;
        RECT 7.000 4.800 7.400 5.200 ;
        RECT 18.200 4.800 18.600 5.200 ;
        RECT 31.800 5.800 32.200 6.200 ;
        RECT 61.400 16.800 61.800 17.200 ;
        RECT 79.000 44.800 79.400 45.200 ;
        RECT 74.200 31.800 74.600 32.200 ;
        RECT 111.000 102.800 111.400 103.200 ;
        RECT 109.400 96.800 109.800 97.200 ;
        RECT 139.000 115.800 139.400 116.200 ;
        RECT 107.000 92.800 107.400 93.200 ;
        RECT 124.600 94.800 125.000 95.200 ;
        RECT 131.000 96.800 131.400 97.200 ;
        RECT 148.600 104.800 149.000 105.200 ;
        RECT 146.200 93.800 146.600 94.200 ;
        RECT 145.400 85.800 145.800 86.200 ;
        RECT 146.200 83.800 146.600 84.200 ;
        RECT 122.200 76.800 122.600 77.200 ;
        RECT 104.600 72.800 105.000 73.200 ;
        RECT 106.200 72.800 106.600 73.200 ;
        RECT 128.600 65.800 129.000 66.200 ;
        RECT 131.800 64.800 132.200 65.200 ;
        RECT 94.200 56.800 94.600 57.200 ;
        RECT 109.400 58.800 109.800 59.200 ;
        RECT 90.200 51.800 90.600 52.200 ;
        RECT 87.000 47.800 87.400 48.200 ;
        RECT 101.400 52.800 101.800 53.200 ;
        RECT 115.000 56.800 115.400 57.200 ;
        RECT 146.200 76.800 146.600 77.200 ;
        RECT 142.200 65.800 142.600 66.200 ;
        RECT 143.000 64.800 143.400 65.200 ;
        RECT 130.200 57.800 130.600 58.200 ;
        RECT 128.600 54.800 129.000 55.200 ;
        RECT 122.200 52.800 122.600 53.200 ;
        RECT 89.400 45.800 89.800 46.200 ;
        RECT 89.400 33.800 89.800 34.200 ;
        RECT 105.400 34.800 105.800 35.200 ;
        RECT 103.000 33.800 103.400 34.200 ;
        RECT 97.400 25.800 97.800 26.200 ;
        RECT 125.400 46.800 125.800 47.200 ;
        RECT 124.600 35.800 125.000 36.200 ;
        RECT 137.400 56.800 137.800 57.200 ;
        RECT 132.600 51.800 133.000 52.200 ;
        RECT 138.200 46.800 138.600 47.200 ;
        RECT 123.000 34.800 123.400 35.200 ;
        RECT 106.200 25.800 106.600 26.200 ;
        RECT 109.400 25.800 109.800 26.200 ;
        RECT 105.400 14.800 105.800 15.200 ;
        RECT 83.000 12.800 83.400 13.200 ;
        RECT 117.400 26.800 117.800 27.200 ;
        RECT 123.800 14.800 124.200 15.200 ;
        RECT 131.800 26.800 132.200 27.200 ;
        RECT 133.400 25.800 133.800 26.200 ;
        RECT 148.600 53.800 149.000 54.200 ;
        RECT 144.600 43.800 145.000 44.200 ;
        RECT 146.200 36.800 146.600 37.200 ;
        RECT 143.800 26.800 144.200 27.200 ;
        RECT 139.000 5.800 139.400 6.200 ;
        RECT 147.800 13.800 148.200 14.200 ;
      LAYER metal3 ;
        RECT 17.400 129.100 17.800 129.200 ;
        RECT 30.200 129.100 30.600 129.200 ;
        RECT 17.400 128.800 30.600 129.100 ;
        RECT 1.400 128.100 1.800 128.200 ;
        RECT 5.400 128.100 5.800 128.200 ;
        RECT 1.400 127.800 5.800 128.100 ;
        RECT 61.400 127.800 61.800 128.200 ;
        RECT 107.000 128.100 107.400 128.200 ;
        RECT 109.400 128.100 109.800 128.200 ;
        RECT 107.000 127.800 109.800 128.100 ;
        RECT 117.400 127.800 117.800 128.200 ;
        RECT 121.400 127.800 121.800 128.200 ;
        RECT 135.800 127.800 136.200 128.200 ;
        RECT 147.800 127.800 148.200 128.200 ;
        RECT 11.000 127.100 11.400 127.200 ;
        RECT 16.600 127.100 17.000 127.200 ;
        RECT 11.000 126.800 17.000 127.100 ;
        RECT 20.600 127.100 21.000 127.200 ;
        RECT 21.400 127.100 21.800 127.200 ;
        RECT 20.600 126.800 21.800 127.100 ;
        RECT 34.200 126.800 34.600 127.200 ;
        RECT 37.400 127.100 37.800 127.200 ;
        RECT 61.400 127.100 61.700 127.800 ;
        RECT 37.400 126.800 61.700 127.100 ;
        RECT 70.200 127.100 70.600 127.200 ;
        RECT 80.600 127.100 81.000 127.200 ;
        RECT 87.000 127.100 87.400 127.200 ;
        RECT 70.200 126.800 87.400 127.100 ;
        RECT 93.400 126.800 93.800 127.200 ;
        RECT 98.200 127.100 98.600 127.200 ;
        RECT 106.200 127.100 106.600 127.200 ;
        RECT 117.400 127.100 117.700 127.800 ;
        RECT 98.200 126.800 117.700 127.100 ;
        RECT 121.400 127.100 121.700 127.800 ;
        RECT 135.000 127.100 135.400 127.200 ;
        RECT 121.400 126.800 135.400 127.100 ;
        RECT 135.800 127.100 136.100 127.800 ;
        RECT 147.800 127.200 148.100 127.800 ;
        RECT 137.400 127.100 137.800 127.200 ;
        RECT 135.800 126.800 137.800 127.100 ;
        RECT 147.800 126.800 148.200 127.200 ;
        RECT 6.200 126.100 6.600 126.200 ;
        RECT 7.000 126.100 7.400 126.200 ;
        RECT 6.200 125.800 7.400 126.100 ;
        RECT 8.600 126.100 9.000 126.200 ;
        RECT 10.200 126.100 10.600 126.200 ;
        RECT 8.600 125.800 10.600 126.100 ;
        RECT 14.200 126.100 14.600 126.200 ;
        RECT 34.200 126.100 34.500 126.800 ;
        RECT 14.200 125.800 34.500 126.100 ;
        RECT 43.000 126.100 43.400 126.200 ;
        RECT 43.000 125.800 44.900 126.100 ;
        RECT 26.200 125.100 26.600 125.200 ;
        RECT 28.600 125.100 29.000 125.200 ;
        RECT 30.200 125.100 30.600 125.200 ;
        RECT 26.200 124.800 30.600 125.100 ;
        RECT 31.000 125.100 31.400 125.200 ;
        RECT 35.000 125.100 35.400 125.200 ;
        RECT 41.400 125.100 41.800 125.200 ;
        RECT 44.600 125.100 44.900 125.800 ;
        RECT 47.800 125.800 48.200 126.200 ;
        RECT 58.200 126.100 58.600 126.200 ;
        RECT 58.200 125.800 63.300 126.100 ;
        RECT 47.800 125.100 48.100 125.800 ;
        RECT 31.000 124.800 44.100 125.100 ;
        RECT 44.600 124.800 48.100 125.100 ;
        RECT 63.000 125.200 63.300 125.800 ;
        RECT 79.000 125.800 79.400 126.200 ;
        RECT 86.200 126.100 86.600 126.200 ;
        RECT 88.600 126.100 89.000 126.200 ;
        RECT 86.200 125.800 89.000 126.100 ;
        RECT 90.200 126.100 90.600 126.200 ;
        RECT 92.600 126.100 93.000 126.200 ;
        RECT 90.200 125.800 93.000 126.100 ;
        RECT 93.400 126.100 93.700 126.800 ;
        RECT 101.400 126.100 101.800 126.200 ;
        RECT 93.400 125.800 101.800 126.100 ;
        RECT 104.600 126.100 105.000 126.200 ;
        RECT 109.400 126.100 109.800 126.200 ;
        RECT 104.600 125.800 109.800 126.100 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 112.600 126.100 113.000 126.200 ;
        RECT 113.400 126.100 113.800 126.200 ;
        RECT 112.600 125.800 113.800 126.100 ;
        RECT 122.200 126.100 122.600 126.200 ;
        RECT 131.800 126.100 132.200 126.200 ;
        RECT 135.000 126.100 135.400 126.200 ;
        RECT 122.200 125.800 135.400 126.100 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 79.000 125.100 79.300 125.800 ;
        RECT 111.800 125.100 112.100 125.800 ;
        RECT 79.000 124.800 112.100 125.100 ;
        RECT 126.200 125.100 126.600 125.200 ;
        RECT 127.000 125.100 127.400 125.200 ;
        RECT 126.200 124.800 127.400 125.100 ;
        RECT 135.000 125.100 135.400 125.200 ;
        RECT 139.000 125.100 139.400 125.200 ;
        RECT 135.000 124.800 139.400 125.100 ;
        RECT 43.800 124.200 44.100 124.800 ;
        RECT 43.800 123.800 44.200 124.200 ;
        RECT 46.200 124.100 46.600 124.200 ;
        RECT 52.600 124.100 53.000 124.200 ;
        RECT 59.800 124.100 60.200 124.200 ;
        RECT 46.200 123.800 60.200 124.100 ;
        RECT 75.800 124.100 76.200 124.200 ;
        RECT 91.800 124.100 92.200 124.200 ;
        RECT 106.200 124.100 106.600 124.200 ;
        RECT 75.800 123.800 106.600 124.100 ;
        RECT 125.400 124.100 125.800 124.200 ;
        RECT 128.600 124.100 129.000 124.200 ;
        RECT 125.400 123.800 129.000 124.100 ;
        RECT 131.000 124.100 131.400 124.200 ;
        RECT 138.200 124.100 138.600 124.200 ;
        RECT 131.000 123.800 138.600 124.100 ;
        RECT 45.400 123.100 45.800 123.200 ;
        RECT 51.000 123.100 51.400 123.200 ;
        RECT 53.400 123.100 53.800 123.200 ;
        RECT 45.400 122.800 53.800 123.100 ;
        RECT 72.600 123.100 73.000 123.200 ;
        RECT 95.800 123.100 96.200 123.200 ;
        RECT 72.600 122.800 96.200 123.100 ;
        RECT 96.600 122.800 97.000 123.200 ;
        RECT 123.800 123.100 124.200 123.200 ;
        RECT 135.000 123.100 135.400 123.200 ;
        RECT 123.800 122.800 135.400 123.100 ;
        RECT 39.800 122.100 40.200 122.200 ;
        RECT 40.600 122.100 41.000 122.200 ;
        RECT 74.200 122.100 74.600 122.200 ;
        RECT 39.800 121.800 41.000 122.100 ;
        RECT 69.400 121.800 74.600 122.100 ;
        RECT 79.000 122.100 79.400 122.200 ;
        RECT 94.200 122.100 94.600 122.200 ;
        RECT 79.000 121.800 94.600 122.100 ;
        RECT 96.600 122.100 96.900 122.800 ;
        RECT 132.600 122.100 133.000 122.200 ;
        RECT 137.400 122.100 137.800 122.200 ;
        RECT 96.600 121.800 137.800 122.100 ;
        RECT 139.800 122.100 140.200 122.200 ;
        RECT 147.000 122.100 147.400 122.200 ;
        RECT 139.800 121.800 147.400 122.100 ;
        RECT 69.400 121.200 69.700 121.800 ;
        RECT 69.400 120.800 69.800 121.200 ;
        RECT 95.800 121.100 96.200 121.200 ;
        RECT 97.400 121.100 97.800 121.200 ;
        RECT 95.800 120.800 97.800 121.100 ;
        RECT 111.000 121.100 111.400 121.200 ;
        RECT 133.400 121.100 133.800 121.200 ;
        RECT 136.600 121.100 137.000 121.200 ;
        RECT 139.800 121.100 140.200 121.200 ;
        RECT 111.000 120.800 140.200 121.100 ;
        RECT 87.800 120.100 88.200 120.200 ;
        RECT 92.600 120.100 93.000 120.200 ;
        RECT 98.200 120.100 98.600 120.200 ;
        RECT 87.800 119.800 98.600 120.100 ;
        RECT 135.000 120.100 135.400 120.200 ;
        RECT 141.400 120.100 141.800 120.200 ;
        RECT 135.000 119.800 141.800 120.100 ;
        RECT 93.400 118.800 93.800 119.200 ;
        RECT 94.200 119.100 94.600 119.200 ;
        RECT 100.600 119.100 101.000 119.200 ;
        RECT 107.000 119.100 107.400 119.200 ;
        RECT 94.200 118.800 107.400 119.100 ;
        RECT 112.600 118.800 113.000 119.200 ;
        RECT 125.400 119.100 125.800 119.200 ;
        RECT 145.400 119.100 145.800 119.200 ;
        RECT 125.400 118.800 145.800 119.100 ;
        RECT 93.400 118.100 93.700 118.800 ;
        RECT 95.000 118.100 95.400 118.200 ;
        RECT 104.600 118.100 105.000 118.200 ;
        RECT 93.400 117.800 105.000 118.100 ;
        RECT 112.600 118.100 112.900 118.800 ;
        RECT 119.000 118.100 119.400 118.200 ;
        RECT 122.200 118.100 122.600 118.200 ;
        RECT 124.600 118.100 125.000 118.200 ;
        RECT 127.800 118.100 128.200 118.200 ;
        RECT 112.600 117.800 128.200 118.100 ;
        RECT 135.800 117.800 136.200 118.200 ;
        RECT 86.200 117.100 86.600 117.200 ;
        RECT 89.400 117.100 89.800 117.200 ;
        RECT 86.200 116.800 89.800 117.100 ;
        RECT 91.000 117.100 91.400 117.200 ;
        RECT 118.200 117.100 118.600 117.200 ;
        RECT 121.400 117.100 121.800 117.200 ;
        RECT 126.200 117.100 126.600 117.200 ;
        RECT 91.000 116.800 126.600 117.100 ;
        RECT 135.800 117.100 136.100 117.800 ;
        RECT 142.200 117.100 142.600 117.200 ;
        RECT 135.800 116.800 142.600 117.100 ;
        RECT 143.800 117.100 144.200 117.200 ;
        RECT 145.400 117.100 145.800 117.200 ;
        RECT 143.800 116.800 145.800 117.100 ;
        RECT 17.400 116.100 17.800 116.200 ;
        RECT 19.800 116.100 20.200 116.200 ;
        RECT 17.400 115.800 20.200 116.100 ;
        RECT 26.200 116.100 26.600 116.200 ;
        RECT 31.800 116.100 32.200 116.200 ;
        RECT 26.200 115.800 32.200 116.100 ;
        RECT 51.800 116.100 52.200 116.200 ;
        RECT 52.600 116.100 53.000 116.200 ;
        RECT 51.800 115.800 53.000 116.100 ;
        RECT 54.200 116.100 54.600 116.200 ;
        RECT 55.000 116.100 55.400 116.200 ;
        RECT 58.200 116.100 58.600 116.200 ;
        RECT 54.200 115.800 58.600 116.100 ;
        RECT 65.400 115.800 65.800 116.200 ;
        RECT 81.400 116.100 81.800 116.200 ;
        RECT 87.800 116.100 88.200 116.200 ;
        RECT 81.400 115.800 88.200 116.100 ;
        RECT 90.200 116.100 90.600 116.200 ;
        RECT 95.800 116.100 96.200 116.200 ;
        RECT 99.000 116.100 99.400 116.200 ;
        RECT 90.200 115.800 99.400 116.100 ;
        RECT 139.000 116.100 139.400 116.200 ;
        RECT 141.400 116.100 141.800 116.200 ;
        RECT 146.200 116.100 146.600 116.200 ;
        RECT 139.000 115.800 146.600 116.100 ;
        RECT 148.600 115.800 149.000 116.200 ;
        RECT 15.800 114.800 16.200 115.200 ;
        RECT 28.600 114.800 29.000 115.200 ;
        RECT 39.800 115.100 40.200 115.200 ;
        RECT 41.400 115.100 41.800 115.200 ;
        RECT 39.800 114.800 41.800 115.100 ;
        RECT 44.600 115.100 45.000 115.200 ;
        RECT 47.800 115.100 48.200 115.200 ;
        RECT 44.600 114.800 48.200 115.100 ;
        RECT 59.800 115.100 60.200 115.200 ;
        RECT 65.400 115.100 65.700 115.800 ;
        RECT 148.600 115.200 148.900 115.800 ;
        RECT 59.800 114.800 65.700 115.100 ;
        RECT 67.800 115.100 68.200 115.200 ;
        RECT 126.200 115.100 126.600 115.200 ;
        RECT 135.000 115.100 135.400 115.200 ;
        RECT 67.800 114.800 135.400 115.100 ;
        RECT 137.400 115.100 137.800 115.200 ;
        RECT 138.200 115.100 138.600 115.200 ;
        RECT 137.400 114.800 138.600 115.100 ;
        RECT 148.600 114.800 149.000 115.200 ;
        RECT 9.400 114.100 9.800 114.200 ;
        RECT 15.800 114.100 16.100 114.800 ;
        RECT 17.400 114.100 17.800 114.200 ;
        RECT 9.400 113.800 17.800 114.100 ;
        RECT 20.600 114.100 21.000 114.200 ;
        RECT 28.600 114.100 28.900 114.800 ;
        RECT 20.600 113.800 28.900 114.100 ;
        RECT 43.000 114.100 43.400 114.200 ;
        RECT 47.000 114.100 47.400 114.200 ;
        RECT 50.200 114.100 50.600 114.200 ;
        RECT 43.000 113.800 50.600 114.100 ;
        RECT 55.000 114.100 55.400 114.200 ;
        RECT 56.600 114.100 57.000 114.200 ;
        RECT 55.000 113.800 57.000 114.100 ;
        RECT 85.400 114.100 85.800 114.200 ;
        RECT 86.200 114.100 86.600 114.200 ;
        RECT 85.400 113.800 86.600 114.100 ;
        RECT 90.200 114.100 90.600 114.200 ;
        RECT 96.600 114.100 97.000 114.200 ;
        RECT 90.200 113.800 97.000 114.100 ;
        RECT 98.200 114.100 98.600 114.200 ;
        RECT 112.600 114.100 113.000 114.200 ;
        RECT 98.200 113.800 113.000 114.100 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 123.800 114.100 124.200 114.200 ;
        RECT 143.800 114.100 144.200 114.200 ;
        RECT 123.800 113.800 144.200 114.100 ;
        RECT 23.000 113.100 23.400 113.200 ;
        RECT 6.200 112.800 23.400 113.100 ;
        RECT 39.800 113.100 40.200 113.200 ;
        RECT 43.800 113.100 44.200 113.200 ;
        RECT 39.800 112.800 44.200 113.100 ;
        RECT 55.800 113.100 56.200 113.200 ;
        RECT 60.600 113.100 61.000 113.200 ;
        RECT 61.400 113.100 61.800 113.200 ;
        RECT 55.800 112.800 61.800 113.100 ;
        RECT 96.600 113.100 96.900 113.800 ;
        RECT 119.800 113.200 120.100 113.800 ;
        RECT 99.800 113.100 100.200 113.200 ;
        RECT 96.600 112.800 100.200 113.100 ;
        RECT 119.800 112.800 120.200 113.200 ;
        RECT 125.400 113.100 125.800 113.200 ;
        RECT 128.600 113.100 129.000 113.200 ;
        RECT 125.400 112.800 129.000 113.100 ;
        RECT 146.200 113.100 146.600 113.200 ;
        RECT 146.200 112.800 147.300 113.100 ;
        RECT 5.400 112.100 5.800 112.200 ;
        RECT 6.200 112.100 6.500 112.800 ;
        RECT 147.000 112.200 147.300 112.800 ;
        RECT 5.400 111.800 6.500 112.100 ;
        RECT 7.000 112.100 7.400 112.200 ;
        RECT 10.200 112.100 10.600 112.200 ;
        RECT 16.600 112.100 17.000 112.200 ;
        RECT 7.000 111.800 17.000 112.100 ;
        RECT 39.000 112.100 39.400 112.200 ;
        RECT 40.600 112.100 41.000 112.200 ;
        RECT 39.000 111.800 41.000 112.100 ;
        RECT 41.400 112.100 41.800 112.200 ;
        RECT 43.000 112.100 43.400 112.200 ;
        RECT 41.400 111.800 43.400 112.100 ;
        RECT 72.600 112.100 73.000 112.200 ;
        RECT 82.200 112.100 82.600 112.200 ;
        RECT 72.600 111.800 82.600 112.100 ;
        RECT 93.400 112.100 93.800 112.200 ;
        RECT 101.400 112.100 101.800 112.200 ;
        RECT 107.000 112.100 107.400 112.200 ;
        RECT 93.400 111.800 107.400 112.100 ;
        RECT 118.200 112.100 118.600 112.200 ;
        RECT 130.200 112.100 130.600 112.200 ;
        RECT 118.200 111.800 130.600 112.100 ;
        RECT 134.200 112.100 134.600 112.200 ;
        RECT 141.400 112.100 141.800 112.200 ;
        RECT 134.200 111.800 141.800 112.100 ;
        RECT 144.600 112.100 145.000 112.200 ;
        RECT 146.200 112.100 146.600 112.200 ;
        RECT 144.600 111.800 146.600 112.100 ;
        RECT 147.000 111.800 147.400 112.200 ;
        RECT 1.400 111.100 1.800 111.200 ;
        RECT 8.600 111.100 9.000 111.200 ;
        RECT 19.000 111.100 19.400 111.200 ;
        RECT 1.400 110.800 19.400 111.100 ;
        RECT 78.200 111.100 78.600 111.200 ;
        RECT 89.400 111.100 89.800 111.200 ;
        RECT 97.400 111.100 97.800 111.200 ;
        RECT 78.200 110.800 97.800 111.100 ;
        RECT 2.200 110.100 2.600 110.200 ;
        RECT 8.600 110.100 9.000 110.200 ;
        RECT 2.200 109.800 9.000 110.100 ;
        RECT 29.400 110.100 29.800 110.200 ;
        RECT 41.400 110.100 41.800 110.200 ;
        RECT 29.400 109.800 41.800 110.100 ;
        RECT 42.200 110.100 42.600 110.200 ;
        RECT 43.800 110.100 44.200 110.200 ;
        RECT 42.200 109.800 44.200 110.100 ;
        RECT 139.800 110.100 140.200 110.200 ;
        RECT 148.600 110.100 149.000 110.200 ;
        RECT 139.800 109.800 149.000 110.100 ;
        RECT 149.400 109.800 149.800 110.200 ;
        RECT 149.400 109.200 149.700 109.800 ;
        RECT 3.800 108.800 4.200 109.200 ;
        RECT 20.600 109.100 21.000 109.200 ;
        RECT 35.800 109.100 36.200 109.200 ;
        RECT 20.600 108.800 36.200 109.100 ;
        RECT 40.600 109.100 41.000 109.200 ;
        RECT 43.800 109.100 44.200 109.200 ;
        RECT 50.200 109.100 50.600 109.200 ;
        RECT 40.600 108.800 50.600 109.100 ;
        RECT 92.600 109.100 93.000 109.200 ;
        RECT 101.400 109.100 101.800 109.200 ;
        RECT 92.600 108.800 101.800 109.100 ;
        RECT 119.800 109.100 120.200 109.200 ;
        RECT 136.600 109.100 137.000 109.200 ;
        RECT 119.800 108.800 137.000 109.100 ;
        RECT 140.600 109.100 141.000 109.200 ;
        RECT 142.200 109.100 142.600 109.200 ;
        RECT 140.600 108.800 142.600 109.100 ;
        RECT 149.400 108.800 149.800 109.200 ;
        RECT 3.800 108.100 4.100 108.800 ;
        RECT 7.000 108.100 7.400 108.200 ;
        RECT 3.800 107.800 7.400 108.100 ;
        RECT 35.000 107.800 35.400 108.200 ;
        RECT 87.800 108.100 88.200 108.200 ;
        RECT 91.800 108.100 92.200 108.200 ;
        RECT 87.800 107.800 92.200 108.100 ;
        RECT 97.400 108.100 97.800 108.200 ;
        RECT 115.000 108.100 115.400 108.200 ;
        RECT 97.400 107.800 115.400 108.100 ;
        RECT 133.400 108.100 133.800 108.200 ;
        RECT 141.400 108.100 141.800 108.200 ;
        RECT 133.400 107.800 141.800 108.100 ;
        RECT 145.400 108.100 145.800 108.200 ;
        RECT 149.400 108.100 149.800 108.200 ;
        RECT 145.400 107.800 149.800 108.100 ;
        RECT 35.000 107.200 35.300 107.800 ;
        RECT 16.600 106.800 17.000 107.200 ;
        RECT 35.000 106.800 35.400 107.200 ;
        RECT 36.600 107.100 37.000 107.200 ;
        RECT 43.000 107.100 43.400 107.200 ;
        RECT 36.600 106.800 43.400 107.100 ;
        RECT 48.600 107.100 49.000 107.200 ;
        RECT 55.000 107.100 55.400 107.200 ;
        RECT 48.600 106.800 55.400 107.100 ;
        RECT 81.400 107.100 81.800 107.200 ;
        RECT 98.200 107.100 98.600 107.200 ;
        RECT 81.400 106.800 98.600 107.100 ;
        RECT 99.000 107.100 99.400 107.200 ;
        RECT 112.600 107.100 113.000 107.200 ;
        RECT 99.000 106.800 113.000 107.100 ;
        RECT 128.600 107.100 129.000 107.200 ;
        RECT 143.000 107.100 143.400 107.200 ;
        RECT 128.600 106.800 143.400 107.100 ;
        RECT 147.800 107.100 148.200 107.200 ;
        RECT 150.200 107.100 150.600 107.200 ;
        RECT 147.800 106.800 150.600 107.100 ;
        RECT 10.200 105.800 10.600 106.200 ;
        RECT 16.600 106.100 16.900 106.800 ;
        RECT 98.200 106.200 98.500 106.800 ;
        RECT 23.000 106.100 23.400 106.200 ;
        RECT 16.600 105.800 23.400 106.100 ;
        RECT 44.600 106.100 45.000 106.200 ;
        RECT 46.200 106.100 46.600 106.200 ;
        RECT 44.600 105.800 46.600 106.100 ;
        RECT 53.400 106.100 53.800 106.200 ;
        RECT 61.400 106.100 61.800 106.200 ;
        RECT 66.200 106.100 66.600 106.200 ;
        RECT 53.400 105.800 58.500 106.100 ;
        RECT 10.200 105.100 10.500 105.800 ;
        RECT 58.200 105.200 58.500 105.800 ;
        RECT 61.400 105.800 66.600 106.100 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 77.400 106.100 77.800 106.200 ;
        RECT 79.800 106.100 80.200 106.200 ;
        RECT 77.400 105.800 80.200 106.100 ;
        RECT 83.800 106.100 84.200 106.200 ;
        RECT 87.000 106.100 87.400 106.200 ;
        RECT 83.800 105.800 87.400 106.100 ;
        RECT 91.000 106.100 91.400 106.200 ;
        RECT 95.000 106.100 95.400 106.200 ;
        RECT 91.000 105.800 95.400 106.100 ;
        RECT 98.200 105.800 98.600 106.200 ;
        RECT 107.000 106.100 107.400 106.200 ;
        RECT 118.200 106.100 118.600 106.200 ;
        RECT 119.800 106.100 120.200 106.200 ;
        RECT 127.800 106.100 128.200 106.200 ;
        RECT 107.000 105.800 128.200 106.100 ;
        RECT 129.400 106.100 129.800 106.200 ;
        RECT 132.600 106.100 133.000 106.200 ;
        RECT 144.600 106.100 145.000 106.200 ;
        RECT 129.400 105.800 133.000 106.100 ;
        RECT 138.200 105.800 145.000 106.100 ;
        RECT 146.200 106.100 146.600 106.200 ;
        RECT 147.000 106.100 147.400 106.200 ;
        RECT 146.200 105.800 147.400 106.100 ;
        RECT 61.400 105.200 61.700 105.800 ;
        RECT 68.600 105.200 68.900 105.800 ;
        RECT 138.200 105.200 138.500 105.800 ;
        RECT 21.400 105.100 21.800 105.200 ;
        RECT 10.200 104.800 21.800 105.100 ;
        RECT 36.600 105.100 37.000 105.200 ;
        RECT 44.600 105.100 45.000 105.200 ;
        RECT 36.600 104.800 45.000 105.100 ;
        RECT 58.200 104.800 58.600 105.200 ;
        RECT 61.400 104.800 61.800 105.200 ;
        RECT 68.600 104.800 69.000 105.200 ;
        RECT 89.400 105.100 89.800 105.200 ;
        RECT 90.200 105.100 90.600 105.200 ;
        RECT 95.800 105.100 96.200 105.200 ;
        RECT 89.400 104.800 96.200 105.100 ;
        RECT 96.600 105.100 97.000 105.200 ;
        RECT 104.600 105.100 105.000 105.200 ;
        RECT 107.000 105.100 107.400 105.200 ;
        RECT 96.600 104.800 107.400 105.100 ;
        RECT 107.800 105.100 108.200 105.200 ;
        RECT 111.800 105.100 112.200 105.200 ;
        RECT 107.800 104.800 112.200 105.100 ;
        RECT 115.000 104.800 115.400 105.200 ;
        RECT 119.000 105.100 119.400 105.200 ;
        RECT 125.400 105.100 125.800 105.200 ;
        RECT 136.600 105.100 137.000 105.200 ;
        RECT 119.000 104.800 137.000 105.100 ;
        RECT 138.200 104.800 138.600 105.200 ;
        RECT 142.200 105.100 142.600 105.200 ;
        RECT 146.200 105.100 146.600 105.200 ;
        RECT 142.200 104.800 146.600 105.100 ;
        RECT 148.600 105.100 149.000 105.200 ;
        RECT 151.000 105.100 151.400 105.200 ;
        RECT 148.600 104.800 151.400 105.100 ;
        RECT 54.200 104.100 54.600 104.200 ;
        RECT 56.600 104.100 57.000 104.200 ;
        RECT 54.200 103.800 57.000 104.100 ;
        RECT 66.200 104.100 66.600 104.200 ;
        RECT 75.000 104.100 75.400 104.200 ;
        RECT 66.200 103.800 75.400 104.100 ;
        RECT 85.400 104.100 85.800 104.200 ;
        RECT 88.600 104.100 89.000 104.200 ;
        RECT 85.400 103.800 89.000 104.100 ;
        RECT 97.400 104.100 97.800 104.200 ;
        RECT 103.000 104.100 103.400 104.200 ;
        RECT 97.400 103.800 103.400 104.100 ;
        RECT 104.600 104.100 105.000 104.200 ;
        RECT 106.200 104.100 106.600 104.200 ;
        RECT 104.600 103.800 106.600 104.100 ;
        RECT 108.600 104.100 109.000 104.200 ;
        RECT 111.000 104.100 111.400 104.200 ;
        RECT 108.600 103.800 111.400 104.100 ;
        RECT 115.000 104.100 115.300 104.800 ;
        RECT 117.400 104.100 117.800 104.200 ;
        RECT 121.400 104.100 121.800 104.200 ;
        RECT 127.000 104.100 127.400 104.200 ;
        RECT 115.000 103.800 127.400 104.100 ;
        RECT 88.600 103.100 89.000 103.200 ;
        RECT 90.200 103.100 90.600 103.200 ;
        RECT 94.200 103.100 94.600 103.200 ;
        RECT 111.000 103.100 111.400 103.200 ;
        RECT 116.600 103.100 117.000 103.200 ;
        RECT 87.800 102.800 94.600 103.100 ;
        RECT 110.200 102.800 117.000 103.100 ;
        RECT 119.800 103.100 120.200 103.200 ;
        RECT 123.000 103.100 123.400 103.200 ;
        RECT 119.800 102.800 123.400 103.100 ;
        RECT 123.800 103.100 124.200 103.200 ;
        RECT 124.600 103.100 125.000 103.200 ;
        RECT 134.200 103.100 134.600 103.200 ;
        RECT 123.800 102.800 134.600 103.100 ;
        RECT 64.600 102.100 65.000 102.200 ;
        RECT 65.400 102.100 65.800 102.200 ;
        RECT 64.600 101.800 65.800 102.100 ;
        RECT 67.000 102.100 67.400 102.200 ;
        RECT 70.200 102.100 70.600 102.200 ;
        RECT 67.000 101.800 70.600 102.100 ;
        RECT 82.200 102.100 82.600 102.200 ;
        RECT 96.600 102.100 97.000 102.200 ;
        RECT 82.200 101.800 97.000 102.100 ;
        RECT 103.800 102.100 104.200 102.200 ;
        RECT 117.400 102.100 117.800 102.200 ;
        RECT 103.800 101.800 117.800 102.100 ;
        RECT 83.000 101.100 83.400 101.200 ;
        RECT 105.400 101.100 105.800 101.200 ;
        RECT 83.000 100.800 105.800 101.100 ;
        RECT 124.600 101.100 125.000 101.200 ;
        RECT 130.200 101.100 130.600 101.200 ;
        RECT 124.600 100.800 130.600 101.100 ;
        RECT 105.400 100.200 105.700 100.800 ;
        RECT 35.800 100.100 36.200 100.200 ;
        RECT 37.400 100.100 37.800 100.200 ;
        RECT 35.800 99.800 37.800 100.100 ;
        RECT 87.000 100.100 87.400 100.200 ;
        RECT 104.600 100.100 105.000 100.200 ;
        RECT 87.000 99.800 105.000 100.100 ;
        RECT 105.400 99.800 105.800 100.200 ;
        RECT 127.800 100.100 128.200 100.200 ;
        RECT 135.000 100.100 135.400 100.200 ;
        RECT 137.400 100.100 137.800 100.200 ;
        RECT 140.600 100.100 141.000 100.200 ;
        RECT 127.800 99.800 141.000 100.100 ;
        RECT 85.400 99.100 85.800 99.200 ;
        RECT 131.800 99.100 132.200 99.200 ;
        RECT 135.800 99.100 136.200 99.200 ;
        RECT 139.000 99.100 139.400 99.200 ;
        RECT 84.600 98.800 139.400 99.100 ;
        RECT 74.200 98.100 74.600 98.200 ;
        RECT 83.800 98.100 84.200 98.200 ;
        RECT 95.800 98.100 96.200 98.200 ;
        RECT 74.200 97.800 96.200 98.100 ;
        RECT 99.800 98.100 100.200 98.200 ;
        RECT 103.000 98.100 103.400 98.200 ;
        RECT 108.600 98.100 109.000 98.200 ;
        RECT 99.800 97.800 109.000 98.100 ;
        RECT 112.600 98.100 113.000 98.200 ;
        RECT 123.800 98.100 124.200 98.200 ;
        RECT 127.000 98.100 127.400 98.200 ;
        RECT 131.000 98.100 131.400 98.200 ;
        RECT 112.600 97.800 131.400 98.100 ;
        RECT 79.800 97.100 80.200 97.200 ;
        RECT 85.400 97.100 85.800 97.200 ;
        RECT 79.000 96.800 85.800 97.100 ;
        RECT 87.000 97.100 87.400 97.200 ;
        RECT 93.400 97.100 93.800 97.200 ;
        RECT 94.200 97.100 94.600 97.200 ;
        RECT 101.400 97.100 101.800 97.200 ;
        RECT 87.000 96.800 101.800 97.100 ;
        RECT 109.400 97.100 109.800 97.200 ;
        RECT 111.800 97.100 112.200 97.200 ;
        RECT 119.000 97.100 119.400 97.200 ;
        RECT 109.400 96.800 119.400 97.100 ;
        RECT 125.400 96.800 125.800 97.200 ;
        RECT 128.600 97.100 129.000 97.200 ;
        RECT 131.000 97.100 131.400 97.200 ;
        RECT 132.600 97.100 133.000 97.200 ;
        RECT 128.600 96.800 133.000 97.100 ;
        RECT 143.800 97.100 144.200 97.200 ;
        RECT 147.000 97.100 147.400 97.200 ;
        RECT 147.800 97.100 148.200 97.200 ;
        RECT 143.800 96.800 148.200 97.100 ;
        RECT 9.400 96.100 9.800 96.200 ;
        RECT 11.000 96.100 11.400 96.200 ;
        RECT 9.400 95.800 11.400 96.100 ;
        RECT 13.400 95.800 13.800 96.200 ;
        RECT 19.800 95.800 20.200 96.200 ;
        RECT 43.800 95.800 44.200 96.200 ;
        RECT 58.200 96.100 58.600 96.200 ;
        RECT 60.600 96.100 61.000 96.200 ;
        RECT 58.200 95.800 61.000 96.100 ;
        RECT 75.000 96.100 75.400 96.200 ;
        RECT 82.200 96.100 82.600 96.200 ;
        RECT 75.000 95.800 82.600 96.100 ;
        RECT 88.600 96.100 89.000 96.200 ;
        RECT 89.400 96.100 89.800 96.200 ;
        RECT 88.600 95.800 89.800 96.100 ;
        RECT 96.600 96.100 97.000 96.200 ;
        RECT 98.200 96.100 98.600 96.200 ;
        RECT 105.400 96.100 105.800 96.200 ;
        RECT 111.800 96.100 112.200 96.200 ;
        RECT 96.600 95.800 112.200 96.100 ;
        RECT 116.600 96.100 117.000 96.200 ;
        RECT 121.400 96.100 121.800 96.200 ;
        RECT 116.600 95.800 121.800 96.100 ;
        RECT 125.400 96.100 125.700 96.800 ;
        RECT 131.000 96.100 131.400 96.200 ;
        RECT 125.400 95.800 131.400 96.100 ;
        RECT 150.200 95.800 150.600 96.200 ;
        RECT 2.200 95.100 2.600 95.200 ;
        RECT 5.400 95.100 5.800 95.200 ;
        RECT 2.200 94.800 5.800 95.100 ;
        RECT 13.400 95.100 13.700 95.800 ;
        RECT 19.800 95.100 20.100 95.800 ;
        RECT 43.800 95.200 44.100 95.800 ;
        RECT 150.200 95.200 150.500 95.800 ;
        RECT 13.400 94.800 20.100 95.100 ;
        RECT 26.200 95.100 26.600 95.200 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 40.600 95.100 41.000 95.200 ;
        RECT 26.200 94.800 41.000 95.100 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 46.200 95.100 46.600 95.200 ;
        RECT 61.400 95.100 61.800 95.200 ;
        RECT 46.200 94.800 61.800 95.100 ;
        RECT 68.600 95.100 69.000 95.200 ;
        RECT 71.000 95.100 71.400 95.200 ;
        RECT 73.400 95.100 73.800 95.200 ;
        RECT 68.600 94.800 73.800 95.100 ;
        RECT 83.800 95.100 84.200 95.200 ;
        RECT 87.800 95.100 88.200 95.200 ;
        RECT 83.800 94.800 88.200 95.100 ;
        RECT 93.400 95.100 93.800 95.200 ;
        RECT 107.000 95.100 107.400 95.200 ;
        RECT 93.400 94.800 107.400 95.100 ;
        RECT 111.800 95.100 112.200 95.200 ;
        RECT 115.000 95.100 115.400 95.200 ;
        RECT 111.800 94.800 115.400 95.100 ;
        RECT 121.400 95.100 121.800 95.200 ;
        RECT 124.600 95.100 125.000 95.200 ;
        RECT 127.000 95.100 127.400 95.200 ;
        RECT 121.400 94.800 127.400 95.100 ;
        RECT 131.000 95.100 131.400 95.200 ;
        RECT 133.400 95.100 133.800 95.200 ;
        RECT 131.000 94.800 133.800 95.100 ;
        RECT 136.600 95.100 137.000 95.200 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 136.600 94.800 139.400 95.100 ;
        RECT 145.400 95.100 145.800 95.200 ;
        RECT 148.600 95.100 149.000 95.200 ;
        RECT 145.400 94.800 149.000 95.100 ;
        RECT 150.200 94.800 150.600 95.200 ;
        RECT 8.600 94.100 9.000 94.400 ;
        RECT 3.000 94.000 9.000 94.100 ;
        RECT 29.400 94.100 29.800 94.200 ;
        RECT 30.200 94.100 30.600 94.200 ;
        RECT 3.000 93.800 8.900 94.000 ;
        RECT 29.400 93.800 30.600 94.100 ;
        RECT 56.600 94.100 57.000 94.200 ;
        RECT 60.600 94.100 61.000 94.200 ;
        RECT 56.600 93.800 61.000 94.100 ;
        RECT 63.800 94.100 64.200 94.200 ;
        RECT 70.200 94.100 70.600 94.200 ;
        RECT 72.600 94.100 73.000 94.200 ;
        RECT 63.800 93.800 73.000 94.100 ;
        RECT 75.000 94.100 75.400 94.200 ;
        RECT 83.000 94.100 83.400 94.200 ;
        RECT 75.000 93.800 83.400 94.100 ;
        RECT 94.200 93.800 94.600 94.200 ;
        RECT 98.200 94.100 98.600 94.200 ;
        RECT 99.000 94.100 99.400 94.200 ;
        RECT 98.200 93.800 99.400 94.100 ;
        RECT 101.400 94.100 101.800 94.200 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 101.400 93.800 103.400 94.100 ;
        RECT 106.200 94.100 106.600 94.200 ;
        RECT 107.000 94.100 107.400 94.200 ;
        RECT 110.200 94.100 110.600 94.200 ;
        RECT 106.200 93.800 110.600 94.100 ;
        RECT 116.600 94.100 117.000 94.200 ;
        RECT 119.000 94.100 119.400 94.200 ;
        RECT 116.600 93.800 119.400 94.100 ;
        RECT 134.200 94.100 134.600 94.200 ;
        RECT 146.200 94.100 146.600 94.200 ;
        RECT 147.000 94.100 147.400 94.200 ;
        RECT 134.200 93.800 143.300 94.100 ;
        RECT 146.200 93.800 147.400 94.100 ;
        RECT 147.800 94.100 148.200 94.200 ;
        RECT 150.200 94.100 150.600 94.200 ;
        RECT 147.800 93.800 150.600 94.100 ;
        RECT 3.000 93.200 3.300 93.800 ;
        RECT 94.200 93.200 94.500 93.800 ;
        RECT 143.000 93.200 143.300 93.800 ;
        RECT 3.000 92.800 3.400 93.200 ;
        RECT 37.400 93.100 37.800 93.200 ;
        RECT 38.200 93.100 38.600 93.200 ;
        RECT 37.400 92.800 38.600 93.100 ;
        RECT 40.600 93.100 41.000 93.200 ;
        RECT 55.000 93.100 55.400 93.200 ;
        RECT 59.000 93.100 59.400 93.200 ;
        RECT 40.600 92.800 59.400 93.100 ;
        RECT 63.800 93.100 64.200 93.200 ;
        RECT 64.600 93.100 65.000 93.200 ;
        RECT 63.800 92.800 65.000 93.100 ;
        RECT 67.800 93.100 68.200 93.200 ;
        RECT 71.800 93.100 72.200 93.200 ;
        RECT 75.800 93.100 76.200 93.200 ;
        RECT 67.800 92.800 76.200 93.100 ;
        RECT 94.200 92.800 94.600 93.200 ;
        RECT 103.800 93.100 104.200 93.200 ;
        RECT 107.000 93.100 107.400 93.200 ;
        RECT 119.800 93.100 120.200 93.200 ;
        RECT 103.800 92.800 120.200 93.100 ;
        RECT 120.600 93.100 121.000 93.200 ;
        RECT 123.000 93.100 123.400 93.200 ;
        RECT 120.600 92.800 123.400 93.100 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 36.600 92.100 37.000 92.200 ;
        RECT 52.600 92.100 53.000 92.200 ;
        RECT 36.600 91.800 53.000 92.100 ;
        RECT 63.000 92.100 63.400 92.200 ;
        RECT 68.600 92.100 69.000 92.200 ;
        RECT 63.000 91.800 69.000 92.100 ;
        RECT 84.600 92.100 85.000 92.200 ;
        RECT 90.200 92.100 90.600 92.200 ;
        RECT 84.600 91.800 90.600 92.100 ;
        RECT 91.800 92.100 92.200 92.200 ;
        RECT 103.800 92.100 104.200 92.200 ;
        RECT 91.800 91.800 104.200 92.100 ;
        RECT 128.600 92.100 129.000 92.200 ;
        RECT 129.400 92.100 129.800 92.200 ;
        RECT 131.800 92.100 132.200 92.200 ;
        RECT 128.600 91.800 132.200 92.100 ;
        RECT 47.800 91.100 48.200 91.200 ;
        RECT 50.200 91.100 50.600 91.200 ;
        RECT 47.800 90.800 50.600 91.100 ;
        RECT 71.800 91.100 72.200 91.200 ;
        RECT 86.200 91.100 86.600 91.200 ;
        RECT 71.800 90.800 86.600 91.100 ;
        RECT 90.200 91.100 90.600 91.200 ;
        RECT 97.400 91.100 97.800 91.200 ;
        RECT 90.200 90.800 97.800 91.100 ;
        RECT 103.800 91.100 104.200 91.200 ;
        RECT 114.200 91.100 114.600 91.200 ;
        RECT 103.800 90.800 114.600 91.100 ;
        RECT 66.200 90.100 66.600 90.200 ;
        RECT 68.600 90.100 69.000 90.200 ;
        RECT 66.200 89.800 69.000 90.100 ;
        RECT 85.400 90.100 85.800 90.200 ;
        RECT 86.200 90.100 86.600 90.200 ;
        RECT 85.400 89.800 86.600 90.100 ;
        RECT 143.800 90.100 144.200 90.200 ;
        RECT 147.800 90.100 148.200 90.200 ;
        RECT 143.800 89.800 148.200 90.100 ;
        RECT 151.000 89.800 151.400 90.200 ;
        RECT 151.000 89.200 151.300 89.800 ;
        RECT 11.000 89.100 11.400 89.200 ;
        RECT 21.400 89.100 21.800 89.200 ;
        RECT 67.800 89.100 68.200 89.200 ;
        RECT 11.000 88.800 21.800 89.100 ;
        RECT 65.400 88.800 68.200 89.100 ;
        RECT 75.800 89.100 76.200 89.200 ;
        RECT 91.800 89.100 92.200 89.200 ;
        RECT 75.800 88.800 92.200 89.100 ;
        RECT 96.600 89.100 97.000 89.200 ;
        RECT 104.600 89.100 105.000 89.200 ;
        RECT 96.600 88.800 105.000 89.100 ;
        RECT 111.000 89.100 111.400 89.200 ;
        RECT 123.800 89.100 124.200 89.200 ;
        RECT 111.000 88.800 124.200 89.100 ;
        RECT 143.000 89.100 143.400 89.200 ;
        RECT 145.400 89.100 145.800 89.200 ;
        RECT 147.800 89.100 148.200 89.200 ;
        RECT 143.000 88.800 148.200 89.100 ;
        RECT 151.000 88.800 151.400 89.200 ;
        RECT 65.400 88.200 65.700 88.800 ;
        RECT 10.200 88.100 10.600 88.200 ;
        RECT 11.800 88.100 12.200 88.200 ;
        RECT 13.400 88.100 13.800 88.200 ;
        RECT 15.800 88.100 16.200 88.200 ;
        RECT 18.200 88.100 18.600 88.200 ;
        RECT 10.200 87.800 13.800 88.100 ;
        RECT 15.000 87.800 18.600 88.100 ;
        RECT 50.200 87.800 50.600 88.200 ;
        RECT 57.400 88.100 57.800 88.200 ;
        RECT 58.200 88.100 58.600 88.200 ;
        RECT 57.400 87.800 58.600 88.100 ;
        RECT 65.400 87.800 65.800 88.200 ;
        RECT 86.200 88.100 86.600 88.200 ;
        RECT 96.600 88.100 97.000 88.200 ;
        RECT 86.200 87.800 97.000 88.100 ;
        RECT 107.000 88.100 107.400 88.200 ;
        RECT 110.200 88.100 110.600 88.200 ;
        RECT 107.000 87.800 110.600 88.100 ;
        RECT 116.600 87.800 117.000 88.200 ;
        RECT 117.400 88.100 117.800 88.200 ;
        RECT 121.400 88.100 121.800 88.200 ;
        RECT 117.400 87.800 121.800 88.100 ;
        RECT 141.400 88.100 141.800 88.200 ;
        RECT 143.800 88.100 144.200 88.200 ;
        RECT 141.400 87.800 144.200 88.100 ;
        RECT 144.600 88.100 145.000 88.200 ;
        RECT 148.600 88.100 149.000 88.200 ;
        RECT 144.600 87.800 149.000 88.100 ;
        RECT 43.000 87.100 43.400 87.200 ;
        RECT 50.200 87.100 50.500 87.800 ;
        RECT 43.000 86.800 50.500 87.100 ;
        RECT 63.800 87.100 64.200 87.200 ;
        RECT 65.400 87.100 65.800 87.200 ;
        RECT 63.800 86.800 65.800 87.100 ;
        RECT 67.800 87.100 68.200 87.200 ;
        RECT 80.600 87.100 81.000 87.200 ;
        RECT 67.800 86.800 81.000 87.100 ;
        RECT 82.200 87.100 82.600 87.200 ;
        RECT 83.000 87.100 83.400 87.200 ;
        RECT 91.000 87.100 91.400 87.200 ;
        RECT 82.200 86.800 91.400 87.100 ;
        RECT 94.200 87.100 94.600 87.200 ;
        RECT 95.800 87.100 96.200 87.200 ;
        RECT 94.200 86.800 96.200 87.100 ;
        RECT 98.200 87.100 98.600 87.200 ;
        RECT 101.400 87.100 101.800 87.200 ;
        RECT 107.000 87.100 107.400 87.200 ;
        RECT 112.600 87.100 113.000 87.200 ;
        RECT 115.000 87.100 115.400 87.200 ;
        RECT 98.200 86.800 115.400 87.100 ;
        RECT 116.600 87.100 116.900 87.800 ;
        RECT 126.200 87.100 126.600 87.200 ;
        RECT 116.600 86.800 126.600 87.100 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 132.600 87.100 133.000 87.200 ;
        RECT 140.600 87.100 141.000 87.200 ;
        RECT 131.800 86.800 133.000 87.100 ;
        RECT 138.200 86.800 141.000 87.100 ;
        RECT 144.600 87.100 145.000 87.200 ;
        RECT 146.200 87.100 146.600 87.200 ;
        RECT 144.600 86.800 146.600 87.100 ;
        RECT 71.800 86.200 72.100 86.800 ;
        RECT 138.200 86.200 138.500 86.800 ;
        RECT 7.800 86.100 8.200 86.200 ;
        RECT 11.800 86.100 12.200 86.200 ;
        RECT 7.800 85.800 12.200 86.100 ;
        RECT 19.000 86.100 19.400 86.200 ;
        RECT 21.400 86.100 21.800 86.200 ;
        RECT 19.000 85.800 21.800 86.100 ;
        RECT 48.600 86.100 49.000 86.200 ;
        RECT 48.600 85.800 52.100 86.100 ;
        RECT 71.800 85.800 72.200 86.200 ;
        RECT 74.200 86.100 74.600 86.200 ;
        RECT 77.400 86.100 77.800 86.200 ;
        RECT 74.200 85.800 77.800 86.100 ;
        RECT 89.400 86.100 89.800 86.200 ;
        RECT 95.800 86.100 96.200 86.200 ;
        RECT 97.400 86.100 97.800 86.200 ;
        RECT 102.200 86.100 102.600 86.200 ;
        RECT 106.200 86.100 106.600 86.200 ;
        RECT 109.400 86.100 109.800 86.200 ;
        RECT 89.400 85.800 109.800 86.100 ;
        RECT 111.000 86.100 111.400 86.200 ;
        RECT 127.000 86.100 127.400 86.200 ;
        RECT 111.000 85.800 127.400 86.100 ;
        RECT 130.200 86.100 130.600 86.200 ;
        RECT 135.000 86.100 135.400 86.200 ;
        RECT 138.200 86.100 138.600 86.200 ;
        RECT 130.200 85.800 138.600 86.100 ;
        RECT 139.000 86.100 139.400 86.200 ;
        RECT 143.000 86.100 143.400 86.200 ;
        RECT 145.400 86.100 145.800 86.200 ;
        RECT 139.000 85.800 145.800 86.100 ;
        RECT 51.800 85.200 52.100 85.800 ;
        RECT 139.000 85.200 139.300 85.800 ;
        RECT 2.200 85.100 2.600 85.200 ;
        RECT 3.000 85.100 3.400 85.200 ;
        RECT 2.200 84.800 3.400 85.100 ;
        RECT 7.800 85.100 8.200 85.200 ;
        RECT 10.200 85.100 10.600 85.200 ;
        RECT 7.800 84.800 10.600 85.100 ;
        RECT 17.400 85.100 17.800 85.200 ;
        RECT 27.800 85.100 28.200 85.200 ;
        RECT 17.400 84.800 28.200 85.100 ;
        RECT 51.800 84.800 52.200 85.200 ;
        RECT 71.000 85.100 71.400 85.200 ;
        RECT 82.200 85.100 82.600 85.200 ;
        RECT 71.000 84.800 82.600 85.100 ;
        RECT 90.200 85.100 90.600 85.200 ;
        RECT 108.600 85.100 109.000 85.200 ;
        RECT 90.200 84.800 109.000 85.100 ;
        RECT 111.000 85.100 111.400 85.200 ;
        RECT 118.200 85.100 118.600 85.200 ;
        RECT 111.000 84.800 118.600 85.100 ;
        RECT 123.800 85.100 124.200 85.200 ;
        RECT 131.000 85.100 131.400 85.200 ;
        RECT 123.800 84.800 131.400 85.100 ;
        RECT 139.000 84.800 139.400 85.200 ;
        RECT 143.800 85.100 144.200 85.200 ;
        RECT 146.200 85.100 146.600 85.200 ;
        RECT 143.800 84.800 146.600 85.100 ;
        RECT 8.600 84.100 9.000 84.200 ;
        RECT 3.000 83.800 9.000 84.100 ;
        RECT 27.000 84.100 27.400 84.200 ;
        RECT 31.000 84.100 31.400 84.200 ;
        RECT 27.000 83.800 31.400 84.100 ;
        RECT 64.600 84.100 65.000 84.200 ;
        RECT 68.600 84.100 69.000 84.200 ;
        RECT 73.400 84.100 73.800 84.200 ;
        RECT 64.600 83.800 73.800 84.100 ;
        RECT 74.200 84.100 74.600 84.200 ;
        RECT 76.600 84.100 77.000 84.200 ;
        RECT 89.400 84.100 89.800 84.200 ;
        RECT 74.200 83.800 89.800 84.100 ;
        RECT 101.400 84.100 101.800 84.200 ;
        RECT 105.400 84.100 105.800 84.200 ;
        RECT 101.400 83.800 105.800 84.100 ;
        RECT 118.200 84.100 118.600 84.200 ;
        RECT 130.200 84.100 130.600 84.200 ;
        RECT 133.400 84.100 133.800 84.200 ;
        RECT 118.200 83.800 133.800 84.100 ;
        RECT 136.600 84.100 137.000 84.200 ;
        RECT 139.800 84.100 140.200 84.200 ;
        RECT 136.600 83.800 140.200 84.100 ;
        RECT 145.400 84.100 145.800 84.200 ;
        RECT 146.200 84.100 146.600 84.200 ;
        RECT 145.400 83.800 146.600 84.100 ;
        RECT 147.000 84.100 147.400 84.200 ;
        RECT 149.400 84.100 149.800 84.200 ;
        RECT 147.000 83.800 149.800 84.100 ;
        RECT 3.000 83.200 3.300 83.800 ;
        RECT 3.000 82.800 3.400 83.200 ;
        RECT 7.000 83.100 7.400 83.200 ;
        RECT 15.800 83.100 16.200 83.200 ;
        RECT 91.800 83.100 92.200 83.200 ;
        RECT 94.200 83.100 94.600 83.200 ;
        RECT 113.400 83.100 113.800 83.200 ;
        RECT 117.400 83.100 117.800 83.200 ;
        RECT 7.000 82.800 16.200 83.100 ;
        RECT 88.600 82.800 117.800 83.100 ;
        RECT 120.600 83.100 121.000 83.200 ;
        RECT 124.600 83.100 125.000 83.200 ;
        RECT 120.600 82.800 125.000 83.100 ;
        RECT 130.200 83.100 130.600 83.200 ;
        RECT 135.000 83.100 135.400 83.200 ;
        RECT 148.600 83.100 149.000 83.200 ;
        RECT 130.200 82.800 149.000 83.100 ;
        RECT 88.600 82.200 88.900 82.800 ;
        RECT 58.200 82.100 58.600 82.200 ;
        RECT 59.000 82.100 59.400 82.200 ;
        RECT 63.800 82.100 64.200 82.200 ;
        RECT 58.200 81.800 64.200 82.100 ;
        RECT 88.600 81.800 89.000 82.200 ;
        RECT 96.600 82.100 97.000 82.200 ;
        RECT 121.400 82.100 121.800 82.200 ;
        RECT 95.800 81.800 121.800 82.100 ;
        RECT 87.000 81.100 87.400 81.200 ;
        RECT 94.200 81.100 94.600 81.200 ;
        RECT 95.000 81.100 95.400 81.200 ;
        RECT 87.000 80.800 95.400 81.100 ;
        RECT 135.800 81.100 136.200 81.200 ;
        RECT 141.400 81.100 141.800 81.200 ;
        RECT 135.800 80.800 141.800 81.100 ;
        RECT 88.600 80.100 89.000 80.200 ;
        RECT 96.600 80.100 97.000 80.200 ;
        RECT 111.800 80.100 112.200 80.200 ;
        RECT 88.600 79.800 112.200 80.100 ;
        RECT 139.000 80.100 139.400 80.200 ;
        RECT 139.800 80.100 140.200 80.200 ;
        RECT 139.000 79.800 140.200 80.100 ;
        RECT 36.600 79.100 37.000 79.200 ;
        RECT 57.400 79.100 57.800 79.200 ;
        RECT 36.600 78.800 57.800 79.100 ;
        RECT 89.400 79.100 89.800 79.200 ;
        RECT 99.000 79.100 99.400 79.200 ;
        RECT 89.400 78.800 99.400 79.100 ;
        RECT 139.000 78.800 139.400 79.200 ;
        RECT 57.400 78.100 57.800 78.200 ;
        RECT 84.600 78.100 85.000 78.200 ;
        RECT 57.400 77.800 85.000 78.100 ;
        RECT 99.800 78.100 100.200 78.200 ;
        RECT 114.200 78.100 114.600 78.200 ;
        RECT 119.000 78.100 119.400 78.200 ;
        RECT 120.600 78.100 121.000 78.200 ;
        RECT 99.800 77.800 121.000 78.100 ;
        RECT 124.600 78.100 125.000 78.200 ;
        RECT 126.200 78.100 126.600 78.200 ;
        RECT 124.600 77.800 126.600 78.100 ;
        RECT 135.000 78.100 135.400 78.200 ;
        RECT 139.000 78.100 139.300 78.800 ;
        RECT 135.000 77.800 139.300 78.100 ;
        RECT 139.800 78.100 140.200 78.200 ;
        RECT 139.800 77.800 145.700 78.100 ;
        RECT 145.400 77.200 145.700 77.800 ;
        RECT 28.600 76.800 29.000 77.200 ;
        RECT 58.200 77.100 58.600 77.200 ;
        RECT 59.000 77.100 59.400 77.200 ;
        RECT 58.200 76.800 59.400 77.100 ;
        RECT 60.600 77.100 61.000 77.200 ;
        RECT 62.200 77.100 62.600 77.200 ;
        RECT 60.600 76.800 62.600 77.100 ;
        RECT 63.800 77.100 64.200 77.200 ;
        RECT 64.600 77.100 65.000 77.200 ;
        RECT 63.800 76.800 65.000 77.100 ;
        RECT 68.600 77.100 69.000 77.200 ;
        RECT 72.600 77.100 73.000 77.200 ;
        RECT 79.000 77.100 79.400 77.200 ;
        RECT 85.400 77.100 85.800 77.200 ;
        RECT 68.600 76.800 85.800 77.100 ;
        RECT 91.800 77.100 92.200 77.200 ;
        RECT 100.600 77.100 101.000 77.200 ;
        RECT 102.200 77.100 102.600 77.200 ;
        RECT 91.800 76.800 102.600 77.100 ;
        RECT 107.800 77.100 108.200 77.200 ;
        RECT 111.800 77.100 112.200 77.200 ;
        RECT 115.000 77.100 115.400 77.200 ;
        RECT 107.800 76.800 115.400 77.100 ;
        RECT 122.200 77.100 122.600 77.200 ;
        RECT 123.800 77.100 124.200 77.200 ;
        RECT 127.800 77.100 128.200 77.200 ;
        RECT 122.200 76.800 128.200 77.100 ;
        RECT 128.600 76.800 129.000 77.200 ;
        RECT 139.000 77.100 139.400 77.200 ;
        RECT 139.800 77.100 140.200 77.200 ;
        RECT 139.000 76.800 140.200 77.100 ;
        RECT 142.200 77.100 142.600 77.200 ;
        RECT 144.600 77.100 145.000 77.200 ;
        RECT 142.200 76.800 145.000 77.100 ;
        RECT 145.400 77.100 145.800 77.200 ;
        RECT 146.200 77.100 146.600 77.200 ;
        RECT 147.800 77.100 148.200 77.200 ;
        RECT 145.400 76.800 148.200 77.100 ;
        RECT 15.000 76.100 15.400 76.200 ;
        RECT 17.400 76.100 17.800 76.200 ;
        RECT 18.200 76.100 18.600 76.200 ;
        RECT 15.000 75.800 18.600 76.100 ;
        RECT 28.600 76.100 28.900 76.800 ;
        RECT 41.400 76.100 41.800 76.200 ;
        RECT 28.600 75.800 41.800 76.100 ;
        RECT 62.200 76.100 62.600 76.200 ;
        RECT 67.800 76.100 68.200 76.200 ;
        RECT 70.200 76.100 70.600 76.200 ;
        RECT 62.200 75.800 70.600 76.100 ;
        RECT 71.800 76.100 72.200 76.200 ;
        RECT 79.800 76.100 80.200 76.200 ;
        RECT 71.800 75.800 80.200 76.100 ;
        RECT 83.800 76.100 84.200 76.200 ;
        RECT 95.800 76.100 96.200 76.200 ;
        RECT 98.200 76.100 98.600 76.200 ;
        RECT 83.800 75.800 98.600 76.100 ;
        RECT 113.400 76.100 113.800 76.200 ;
        RECT 116.600 76.100 117.000 76.200 ;
        RECT 113.400 75.800 117.000 76.100 ;
        RECT 127.000 75.800 127.400 76.200 ;
        RECT 128.600 76.100 128.900 76.800 ;
        RECT 131.000 76.100 131.400 76.200 ;
        RECT 128.600 75.800 131.400 76.100 ;
        RECT 138.200 76.100 138.600 76.200 ;
        RECT 140.600 76.100 141.000 76.200 ;
        RECT 143.800 76.100 144.200 76.200 ;
        RECT 138.200 75.800 144.200 76.100 ;
        RECT 147.800 76.100 148.200 76.200 ;
        RECT 149.400 76.100 149.800 76.200 ;
        RECT 147.800 75.800 149.800 76.100 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 3.800 74.800 5.000 75.100 ;
        RECT 34.200 75.100 34.600 75.200 ;
        RECT 43.000 75.100 43.400 75.200 ;
        RECT 34.200 74.800 43.400 75.100 ;
        RECT 59.000 75.100 59.400 75.200 ;
        RECT 64.600 75.100 65.000 75.200 ;
        RECT 67.000 75.100 67.400 75.200 ;
        RECT 71.000 75.100 71.400 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 79.800 75.100 80.200 75.200 ;
        RECT 59.000 74.800 71.400 75.100 ;
        RECT 74.200 74.800 80.200 75.100 ;
        RECT 85.400 75.100 85.800 75.200 ;
        RECT 91.800 75.100 92.200 75.200 ;
        RECT 85.400 74.800 92.200 75.100 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 107.800 75.100 108.200 75.200 ;
        RECT 111.000 75.100 111.400 75.200 ;
        RECT 107.800 74.800 111.400 75.100 ;
        RECT 112.600 75.100 113.000 75.200 ;
        RECT 122.200 75.100 122.600 75.200 ;
        RECT 127.000 75.100 127.300 75.800 ;
        RECT 112.600 74.800 127.300 75.100 ;
        RECT 138.200 75.100 138.600 75.200 ;
        RECT 139.000 75.100 139.400 75.200 ;
        RECT 138.200 74.800 139.400 75.100 ;
        RECT 139.800 75.100 140.200 75.200 ;
        RECT 145.400 75.100 145.800 75.200 ;
        RECT 139.800 74.800 145.800 75.100 ;
        RECT 148.600 74.800 149.000 75.200 ;
        RECT 93.400 74.200 93.700 74.800 ;
        RECT 120.600 74.200 120.900 74.800 ;
        RECT 16.600 73.800 17.000 74.200 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 37.400 74.100 37.800 74.200 ;
        RECT 52.600 74.100 53.000 74.200 ;
        RECT 37.400 73.800 53.000 74.100 ;
        RECT 63.800 74.100 64.200 74.200 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 63.800 73.800 66.600 74.100 ;
        RECT 79.000 74.100 79.400 74.200 ;
        RECT 86.200 74.100 86.600 74.200 ;
        RECT 79.000 73.800 86.600 74.100 ;
        RECT 87.000 74.100 87.400 74.200 ;
        RECT 89.400 74.100 89.800 74.200 ;
        RECT 87.000 73.800 89.800 74.100 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 93.400 73.800 93.800 74.200 ;
        RECT 99.000 74.100 99.400 74.200 ;
        RECT 107.000 74.100 107.400 74.200 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 99.000 73.800 109.000 74.100 ;
        RECT 120.600 73.800 121.000 74.200 ;
        RECT 124.600 74.100 125.000 74.200 ;
        RECT 128.600 74.100 129.000 74.200 ;
        RECT 124.600 73.800 129.000 74.100 ;
        RECT 137.400 73.800 137.800 74.200 ;
        RECT 147.000 74.100 147.400 74.200 ;
        RECT 148.600 74.100 148.900 74.800 ;
        RECT 147.000 73.800 148.900 74.100 ;
        RECT 150.200 73.800 150.600 74.200 ;
        RECT 12.600 73.100 13.000 73.200 ;
        RECT 16.600 73.100 16.900 73.800 ;
        RECT 12.600 72.800 16.900 73.100 ;
        RECT 20.600 73.200 20.900 73.800 ;
        RECT 90.200 73.200 90.500 73.800 ;
        RECT 137.400 73.200 137.700 73.800 ;
        RECT 150.200 73.200 150.500 73.800 ;
        RECT 20.600 72.800 21.000 73.200 ;
        RECT 63.000 73.100 63.400 73.200 ;
        RECT 64.600 73.100 65.000 73.200 ;
        RECT 63.000 72.800 65.000 73.100 ;
        RECT 90.200 72.800 90.600 73.200 ;
        RECT 91.000 73.100 91.400 73.200 ;
        RECT 98.200 73.100 98.600 73.200 ;
        RECT 91.000 72.800 98.600 73.100 ;
        RECT 104.600 73.100 105.000 73.200 ;
        RECT 106.200 73.100 106.600 73.200 ;
        RECT 111.000 73.100 111.400 73.200 ;
        RECT 104.600 72.800 111.400 73.100 ;
        RECT 112.600 73.100 113.000 73.200 ;
        RECT 119.800 73.100 120.200 73.200 ;
        RECT 112.600 72.800 120.200 73.100 ;
        RECT 120.600 73.100 121.000 73.200 ;
        RECT 124.600 73.100 125.000 73.200 ;
        RECT 126.200 73.100 126.600 73.200 ;
        RECT 120.600 72.800 126.600 73.100 ;
        RECT 137.400 72.800 137.800 73.200 ;
        RECT 150.200 72.800 150.600 73.200 ;
        RECT 2.200 72.100 2.600 72.200 ;
        RECT 3.800 72.100 4.200 72.200 ;
        RECT 1.400 71.800 4.200 72.100 ;
        RECT 48.600 72.100 49.000 72.200 ;
        RECT 59.000 72.100 59.400 72.200 ;
        RECT 48.600 71.800 59.400 72.100 ;
        RECT 59.800 72.100 60.200 72.200 ;
        RECT 87.800 72.100 88.200 72.200 ;
        RECT 101.400 72.100 101.800 72.200 ;
        RECT 59.800 71.800 88.200 72.100 ;
        RECT 94.200 71.800 101.800 72.100 ;
        RECT 21.400 71.100 21.800 71.200 ;
        RECT 30.200 71.100 30.600 71.200 ;
        RECT 21.400 70.800 30.600 71.100 ;
        RECT 35.800 71.100 36.200 71.200 ;
        RECT 40.600 71.100 41.000 71.200 ;
        RECT 35.800 70.800 41.000 71.100 ;
        RECT 59.000 71.100 59.400 71.200 ;
        RECT 73.400 71.100 73.800 71.200 ;
        RECT 59.000 70.800 73.800 71.100 ;
        RECT 82.200 71.100 82.600 71.200 ;
        RECT 94.200 71.100 94.500 71.800 ;
        RECT 82.200 70.800 94.500 71.100 ;
        RECT 17.400 69.800 17.800 70.200 ;
        RECT 84.600 70.100 85.000 70.200 ;
        RECT 91.000 70.100 91.400 70.200 ;
        RECT 84.600 69.800 91.400 70.100 ;
        RECT 17.400 69.200 17.700 69.800 ;
        RECT 4.600 69.100 5.000 69.200 ;
        RECT 12.600 69.100 13.000 69.200 ;
        RECT 4.600 68.800 13.000 69.100 ;
        RECT 17.400 68.800 17.800 69.200 ;
        RECT 32.600 69.100 33.000 69.200 ;
        RECT 39.800 69.100 40.200 69.200 ;
        RECT 32.600 68.800 40.200 69.100 ;
        RECT 58.200 69.100 58.600 69.200 ;
        RECT 60.600 69.100 61.000 69.200 ;
        RECT 58.200 68.800 61.000 69.100 ;
        RECT 93.400 68.800 93.800 69.200 ;
        RECT 99.000 69.100 99.400 69.200 ;
        RECT 103.000 69.100 103.400 69.200 ;
        RECT 99.000 68.800 103.400 69.100 ;
        RECT 119.800 69.100 120.200 69.200 ;
        RECT 126.200 69.100 126.600 69.200 ;
        RECT 119.800 68.800 126.600 69.100 ;
        RECT 143.000 69.100 143.400 69.200 ;
        RECT 146.200 69.100 146.600 69.200 ;
        RECT 143.000 68.800 146.600 69.100 ;
        RECT 9.400 68.100 9.800 68.200 ;
        RECT 17.400 68.100 17.800 68.200 ;
        RECT 9.400 67.800 17.800 68.100 ;
        RECT 28.600 67.800 29.000 68.200 ;
        RECT 49.400 67.800 49.800 68.200 ;
        RECT 66.200 68.100 66.600 68.200 ;
        RECT 73.400 68.100 73.800 68.200 ;
        RECT 66.200 67.800 73.800 68.100 ;
        RECT 76.600 68.100 77.000 68.200 ;
        RECT 77.400 68.100 77.800 68.200 ;
        RECT 76.600 67.800 77.800 68.100 ;
        RECT 83.800 68.100 84.200 68.200 ;
        RECT 85.400 68.100 85.800 68.200 ;
        RECT 91.000 68.100 91.400 68.200 ;
        RECT 83.800 67.800 91.400 68.100 ;
        RECT 91.800 67.800 92.200 68.200 ;
        RECT 93.400 68.100 93.700 68.800 ;
        RECT 107.800 68.100 108.200 68.200 ;
        RECT 112.600 68.100 113.000 68.200 ;
        RECT 93.400 67.800 107.300 68.100 ;
        RECT 107.800 67.800 113.000 68.100 ;
        RECT 115.000 68.100 115.400 68.200 ;
        RECT 119.000 68.100 119.400 68.200 ;
        RECT 121.400 68.100 121.800 68.200 ;
        RECT 115.000 67.800 121.800 68.100 ;
        RECT 124.600 67.800 125.000 68.200 ;
        RECT 138.200 68.100 138.600 68.200 ;
        RECT 125.400 67.800 138.600 68.100 ;
        RECT 146.200 67.800 146.600 68.200 ;
        RECT 2.200 67.100 2.600 67.200 ;
        RECT 8.600 67.100 9.000 67.200 ;
        RECT 2.200 66.800 9.000 67.100 ;
        RECT 10.200 67.100 10.600 67.200 ;
        RECT 11.000 67.100 11.400 67.200 ;
        RECT 28.600 67.100 28.900 67.800 ;
        RECT 10.200 66.800 28.900 67.100 ;
        RECT 43.000 67.100 43.400 67.200 ;
        RECT 49.400 67.100 49.700 67.800 ;
        RECT 91.800 67.200 92.100 67.800 ;
        RECT 43.000 66.800 49.700 67.100 ;
        RECT 63.800 67.100 64.200 67.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 67.800 67.100 68.200 67.200 ;
        RECT 63.800 66.800 68.200 67.100 ;
        RECT 68.600 67.100 69.000 67.200 ;
        RECT 79.000 67.100 79.400 67.200 ;
        RECT 68.600 66.800 79.400 67.100 ;
        RECT 88.600 67.100 89.000 67.200 ;
        RECT 89.400 67.100 89.800 67.200 ;
        RECT 88.600 66.800 89.800 67.100 ;
        RECT 91.800 66.800 92.200 67.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 106.200 67.100 106.600 67.200 ;
        RECT 94.200 66.800 106.600 67.100 ;
        RECT 107.000 67.100 107.300 67.800 ;
        RECT 124.600 67.200 124.900 67.800 ;
        RECT 125.400 67.200 125.700 67.800 ;
        RECT 120.600 67.100 121.000 67.200 ;
        RECT 107.000 66.800 121.000 67.100 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 122.200 67.100 122.600 67.200 ;
        RECT 124.600 67.100 125.000 67.200 ;
        RECT 122.200 66.800 125.000 67.100 ;
        RECT 125.400 66.800 125.800 67.200 ;
        RECT 137.400 67.100 137.800 67.200 ;
        RECT 146.200 67.100 146.500 67.800 ;
        RECT 137.400 66.800 146.500 67.100 ;
        RECT 8.600 66.100 8.900 66.800 ;
        RECT 15.000 66.100 15.400 66.200 ;
        RECT 8.600 65.800 15.400 66.100 ;
        RECT 15.800 66.100 16.200 66.200 ;
        RECT 23.800 66.100 24.200 66.200 ;
        RECT 15.800 65.800 24.200 66.100 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 62.200 66.100 62.600 66.200 ;
        RECT 65.400 66.100 65.800 66.200 ;
        RECT 69.400 66.100 69.800 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 31.800 65.800 51.300 66.100 ;
        RECT 62.200 65.800 77.000 66.100 ;
        RECT 79.800 66.100 80.200 66.200 ;
        RECT 99.800 66.100 100.200 66.200 ;
        RECT 79.800 65.800 100.200 66.100 ;
        RECT 103.800 66.100 104.200 66.200 ;
        RECT 110.200 66.100 110.600 66.200 ;
        RECT 103.800 65.800 110.600 66.100 ;
        RECT 115.800 66.100 116.200 66.200 ;
        RECT 121.400 66.100 121.700 66.800 ;
        RECT 123.000 66.100 123.400 66.200 ;
        RECT 128.600 66.100 129.000 66.200 ;
        RECT 115.800 65.800 129.000 66.100 ;
        RECT 131.000 66.100 131.400 66.200 ;
        RECT 133.400 66.100 133.800 66.200 ;
        RECT 131.000 65.800 133.800 66.100 ;
        RECT 142.200 66.100 142.600 66.200 ;
        RECT 143.800 66.100 144.200 66.200 ;
        RECT 142.200 65.800 144.200 66.100 ;
        RECT 51.000 65.200 51.300 65.800 ;
        RECT 15.000 65.100 15.400 65.200 ;
        RECT 15.800 65.100 16.200 65.200 ;
        RECT 23.000 65.100 23.400 65.200 ;
        RECT 15.000 64.800 23.400 65.100 ;
        RECT 51.000 64.800 51.400 65.200 ;
        RECT 60.600 65.100 61.000 65.200 ;
        RECT 61.400 65.100 61.800 65.200 ;
        RECT 60.600 64.800 61.800 65.100 ;
        RECT 64.600 65.100 65.000 65.200 ;
        RECT 76.600 65.100 77.000 65.200 ;
        RECT 64.600 64.800 77.000 65.100 ;
        RECT 77.400 65.100 77.800 65.200 ;
        RECT 80.600 65.100 81.000 65.200 ;
        RECT 77.400 64.800 81.000 65.100 ;
        RECT 90.200 65.100 90.600 65.200 ;
        RECT 93.400 65.100 93.800 65.200 ;
        RECT 103.000 65.100 103.400 65.200 ;
        RECT 90.200 64.800 103.400 65.100 ;
        RECT 115.800 65.100 116.200 65.200 ;
        RECT 117.400 65.100 117.800 65.200 ;
        RECT 119.000 65.100 119.400 65.200 ;
        RECT 119.800 65.100 120.200 65.200 ;
        RECT 115.800 64.800 118.500 65.100 ;
        RECT 119.000 64.800 120.200 65.100 ;
        RECT 124.600 65.100 125.000 65.200 ;
        RECT 128.600 65.100 129.000 65.200 ;
        RECT 124.600 64.800 129.000 65.100 ;
        RECT 129.400 65.100 129.800 65.200 ;
        RECT 130.200 65.100 130.600 65.200 ;
        RECT 129.400 64.800 130.600 65.100 ;
        RECT 131.800 65.100 132.200 65.200 ;
        RECT 135.000 65.100 135.400 65.200 ;
        RECT 137.400 65.100 137.800 65.200 ;
        RECT 131.800 64.800 137.800 65.100 ;
        RECT 143.000 65.100 143.400 65.200 ;
        RECT 145.400 65.100 145.800 65.200 ;
        RECT 143.000 64.800 145.800 65.100 ;
        RECT 19.000 64.100 19.400 64.200 ;
        RECT 29.400 64.100 29.800 64.200 ;
        RECT 19.000 63.800 29.800 64.100 ;
        RECT 71.800 64.100 72.200 64.200 ;
        RECT 79.000 64.100 79.400 64.200 ;
        RECT 71.800 63.800 79.400 64.100 ;
        RECT 80.600 64.100 81.000 64.200 ;
        RECT 114.200 64.100 114.600 64.200 ;
        RECT 133.400 64.100 133.800 64.200 ;
        RECT 136.600 64.100 137.000 64.200 ;
        RECT 80.600 63.800 137.000 64.100 ;
        RECT 47.800 63.100 48.200 63.200 ;
        RECT 70.200 63.100 70.600 63.200 ;
        RECT 79.800 63.100 80.200 63.200 ;
        RECT 88.600 63.100 89.000 63.200 ;
        RECT 47.800 62.800 89.000 63.100 ;
        RECT 133.400 63.100 133.800 63.200 ;
        RECT 140.600 63.100 141.000 63.200 ;
        RECT 133.400 62.800 141.000 63.100 ;
        RECT 55.000 62.100 55.400 62.200 ;
        RECT 63.800 62.100 64.200 62.200 ;
        RECT 67.000 62.100 67.400 62.200 ;
        RECT 55.000 61.800 67.400 62.100 ;
        RECT 77.400 62.100 77.800 62.200 ;
        RECT 96.600 62.100 97.000 62.200 ;
        RECT 77.400 61.800 97.000 62.100 ;
        RECT 52.600 61.100 53.000 61.200 ;
        RECT 72.600 61.100 73.000 61.200 ;
        RECT 52.600 60.800 73.000 61.100 ;
        RECT 98.200 61.100 98.600 61.200 ;
        RECT 108.600 61.100 109.000 61.200 ;
        RECT 98.200 60.800 109.000 61.100 ;
        RECT 51.000 60.100 51.400 60.200 ;
        RECT 58.200 60.100 58.600 60.200 ;
        RECT 51.000 59.800 58.600 60.100 ;
        RECT 70.200 60.100 70.600 60.200 ;
        RECT 132.600 60.100 133.000 60.200 ;
        RECT 139.800 60.100 140.200 60.200 ;
        RECT 151.000 60.100 151.400 60.200 ;
        RECT 70.200 59.800 151.400 60.100 ;
        RECT 11.000 59.100 11.400 59.200 ;
        RECT 12.600 59.100 13.000 59.200 ;
        RECT 31.800 59.100 32.200 59.200 ;
        RECT 55.800 59.100 56.200 59.200 ;
        RECT 11.000 58.800 13.000 59.100 ;
        RECT 31.000 58.800 56.200 59.100 ;
        RECT 91.000 59.100 91.400 59.200 ;
        RECT 92.600 59.100 93.000 59.200 ;
        RECT 106.200 59.100 106.600 59.200 ;
        RECT 91.000 58.800 106.600 59.100 ;
        RECT 109.400 59.100 109.800 59.200 ;
        RECT 112.600 59.100 113.000 59.200 ;
        RECT 131.000 59.100 131.400 59.200 ;
        RECT 109.400 58.800 131.400 59.100 ;
        RECT 143.000 59.100 143.400 59.200 ;
        RECT 147.000 59.100 147.400 59.200 ;
        RECT 143.000 58.800 147.400 59.100 ;
        RECT 47.800 58.100 48.200 58.200 ;
        RECT 54.200 58.100 54.600 58.200 ;
        RECT 47.800 57.800 54.600 58.100 ;
        RECT 103.800 57.800 104.200 58.200 ;
        RECT 107.800 58.100 108.200 58.200 ;
        RECT 110.200 58.100 110.600 58.200 ;
        RECT 113.400 58.100 113.800 58.200 ;
        RECT 115.000 58.100 115.400 58.200 ;
        RECT 107.800 57.800 115.400 58.100 ;
        RECT 123.800 58.100 124.200 58.200 ;
        RECT 130.200 58.100 130.600 58.200 ;
        RECT 135.800 58.100 136.200 58.200 ;
        RECT 144.600 58.100 145.000 58.200 ;
        RECT 123.800 57.800 128.900 58.100 ;
        RECT 129.400 57.800 145.000 58.100 ;
        RECT 148.600 57.800 149.000 58.200 ;
        RECT 24.600 56.800 25.000 57.200 ;
        RECT 50.200 57.100 50.600 57.200 ;
        RECT 55.800 57.100 56.200 57.200 ;
        RECT 59.000 57.100 59.400 57.200 ;
        RECT 61.400 57.100 61.800 57.200 ;
        RECT 50.200 56.800 61.800 57.100 ;
        RECT 63.000 56.800 63.400 57.200 ;
        RECT 65.400 57.100 65.800 57.200 ;
        RECT 66.200 57.100 66.600 57.200 ;
        RECT 74.200 57.100 74.600 57.200 ;
        RECT 65.400 56.800 74.600 57.100 ;
        RECT 90.200 57.100 90.600 57.200 ;
        RECT 94.200 57.100 94.600 57.200 ;
        RECT 99.000 57.100 99.400 57.200 ;
        RECT 90.200 56.800 99.400 57.100 ;
        RECT 103.800 57.100 104.100 57.800 ;
        RECT 106.200 57.100 106.600 57.200 ;
        RECT 103.800 56.800 106.600 57.100 ;
        RECT 111.800 57.100 112.200 57.200 ;
        RECT 115.000 57.100 115.400 57.200 ;
        RECT 116.600 57.100 117.000 57.200 ;
        RECT 111.800 56.800 117.000 57.100 ;
        RECT 118.200 57.100 118.600 57.200 ;
        RECT 124.600 57.100 125.000 57.200 ;
        RECT 127.800 57.100 128.200 57.200 ;
        RECT 118.200 56.800 128.200 57.100 ;
        RECT 128.600 57.100 128.900 57.800 ;
        RECT 131.000 57.100 131.400 57.200 ;
        RECT 128.600 56.800 131.400 57.100 ;
        RECT 135.000 56.800 135.400 57.200 ;
        RECT 137.400 57.100 137.800 57.200 ;
        RECT 148.600 57.100 148.900 57.800 ;
        RECT 137.400 56.800 148.900 57.100 ;
        RECT 3.800 55.800 4.200 56.200 ;
        RECT 8.600 55.800 9.000 56.200 ;
        RECT 24.600 56.100 24.900 56.800 ;
        RECT 29.400 56.100 29.800 56.200 ;
        RECT 35.000 56.100 35.400 56.200 ;
        RECT 24.600 55.800 35.400 56.100 ;
        RECT 52.600 56.100 53.000 56.200 ;
        RECT 54.200 56.100 54.600 56.200 ;
        RECT 52.600 55.800 54.600 56.100 ;
        RECT 59.000 56.100 59.400 56.200 ;
        RECT 63.000 56.100 63.300 56.800 ;
        RECT 135.000 56.200 135.300 56.800 ;
        RECT 74.200 56.100 74.600 56.200 ;
        RECT 104.600 56.100 105.000 56.200 ;
        RECT 59.000 55.800 74.600 56.100 ;
        RECT 94.200 55.800 105.000 56.100 ;
        RECT 107.000 56.100 107.400 56.200 ;
        RECT 123.000 56.100 123.400 56.200 ;
        RECT 125.400 56.100 125.800 56.200 ;
        RECT 107.000 55.800 125.800 56.100 ;
        RECT 135.000 55.800 135.400 56.200 ;
        RECT 147.800 55.800 148.200 56.200 ;
        RECT 3.800 55.100 4.100 55.800 ;
        RECT 8.600 55.100 8.900 55.800 ;
        RECT 94.200 55.200 94.500 55.800 ;
        RECT 147.800 55.200 148.100 55.800 ;
        RECT 3.800 54.800 8.900 55.100 ;
        RECT 23.800 55.100 24.200 55.200 ;
        RECT 26.200 55.100 26.600 55.200 ;
        RECT 27.800 55.100 28.200 55.200 ;
        RECT 23.800 54.800 28.200 55.100 ;
        RECT 39.800 54.800 40.200 55.200 ;
        RECT 51.000 55.100 51.400 55.200 ;
        RECT 54.200 55.100 54.600 55.200 ;
        RECT 51.000 54.800 54.600 55.100 ;
        RECT 60.600 55.100 61.000 55.200 ;
        RECT 63.800 55.100 64.200 55.200 ;
        RECT 60.600 54.800 64.200 55.100 ;
        RECT 68.600 55.100 69.000 55.200 ;
        RECT 77.400 55.100 77.800 55.200 ;
        RECT 68.600 54.800 77.800 55.100 ;
        RECT 87.000 55.100 87.400 55.200 ;
        RECT 88.600 55.100 89.000 55.200 ;
        RECT 87.000 54.800 89.000 55.100 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 95.800 55.100 96.200 55.200 ;
        RECT 99.000 55.100 99.400 55.200 ;
        RECT 95.800 54.800 99.400 55.100 ;
        RECT 101.400 55.100 101.800 55.200 ;
        RECT 114.200 55.100 114.600 55.200 ;
        RECT 101.400 54.800 114.600 55.100 ;
        RECT 117.400 55.100 117.800 55.200 ;
        RECT 123.000 55.100 123.400 55.200 ;
        RECT 127.000 55.100 127.400 55.200 ;
        RECT 117.400 54.800 127.400 55.100 ;
        RECT 128.600 55.100 129.000 55.200 ;
        RECT 134.200 55.100 134.600 55.200 ;
        RECT 128.600 54.800 134.600 55.100 ;
        RECT 147.800 55.100 148.200 55.200 ;
        RECT 149.400 55.100 149.800 55.200 ;
        RECT 147.800 54.800 149.800 55.100 ;
        RECT 32.600 54.100 33.000 54.200 ;
        RECT 39.800 54.100 40.100 54.800 ;
        RECT 32.600 53.800 40.100 54.100 ;
        RECT 42.200 54.100 42.600 54.200 ;
        RECT 53.400 54.100 53.800 54.200 ;
        RECT 42.200 53.800 53.800 54.100 ;
        RECT 56.600 54.100 57.000 54.200 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 59.000 54.100 59.400 54.200 ;
        RECT 56.600 53.800 59.400 54.100 ;
        RECT 62.200 54.100 62.600 54.200 ;
        RECT 65.400 54.100 65.800 54.200 ;
        RECT 62.200 53.800 65.800 54.100 ;
        RECT 75.000 54.100 75.400 54.200 ;
        RECT 87.000 54.100 87.400 54.200 ;
        RECT 75.000 53.800 87.400 54.100 ;
        RECT 87.800 54.100 88.200 54.200 ;
        RECT 97.400 54.100 97.800 54.200 ;
        RECT 87.800 53.800 97.800 54.100 ;
        RECT 98.200 54.100 98.600 54.200 ;
        RECT 101.400 54.100 101.800 54.200 ;
        RECT 98.200 53.800 101.800 54.100 ;
        RECT 102.200 54.100 102.600 54.200 ;
        RECT 103.000 54.100 103.400 54.200 ;
        RECT 102.200 53.800 103.400 54.100 ;
        RECT 117.400 54.100 117.800 54.200 ;
        RECT 119.000 54.100 119.400 54.200 ;
        RECT 129.400 54.100 129.800 54.200 ;
        RECT 117.400 53.800 119.400 54.100 ;
        RECT 123.000 53.800 129.800 54.100 ;
        RECT 139.800 54.100 140.200 54.200 ;
        RECT 140.600 54.100 141.000 54.200 ;
        RECT 139.800 53.800 141.000 54.100 ;
        RECT 146.200 54.100 146.600 54.200 ;
        RECT 148.600 54.100 149.000 54.200 ;
        RECT 146.200 53.800 149.000 54.100 ;
        RECT 123.000 53.200 123.300 53.800 ;
        RECT 3.000 53.100 3.400 53.200 ;
        RECT 8.600 53.100 9.000 53.200 ;
        RECT 3.000 52.800 9.000 53.100 ;
        RECT 15.000 53.100 15.400 53.200 ;
        RECT 17.400 53.100 17.800 53.200 ;
        RECT 15.000 52.800 17.800 53.100 ;
        RECT 21.400 53.100 21.800 53.200 ;
        RECT 24.600 53.100 25.000 53.200 ;
        RECT 26.200 53.100 26.600 53.200 ;
        RECT 21.400 52.800 26.600 53.100 ;
        RECT 63.000 53.100 63.400 53.200 ;
        RECT 66.200 53.100 66.600 53.200 ;
        RECT 63.000 52.800 66.600 53.100 ;
        RECT 79.800 53.100 80.200 53.200 ;
        RECT 80.600 53.100 81.000 53.200 ;
        RECT 81.400 53.100 81.800 53.200 ;
        RECT 87.800 53.100 88.200 53.200 ;
        RECT 91.800 53.100 92.200 53.200 ;
        RECT 79.800 52.800 81.800 53.100 ;
        RECT 87.000 52.800 92.200 53.100 ;
        RECT 96.600 53.100 97.000 53.200 ;
        RECT 101.400 53.100 101.800 53.200 ;
        RECT 103.800 53.100 104.200 53.200 ;
        RECT 96.600 52.800 104.200 53.100 ;
        RECT 107.800 53.100 108.200 53.200 ;
        RECT 119.800 53.100 120.200 53.200 ;
        RECT 107.800 52.800 120.200 53.100 ;
        RECT 122.200 53.100 122.600 53.200 ;
        RECT 123.000 53.100 123.400 53.200 ;
        RECT 127.800 53.100 128.200 53.200 ;
        RECT 128.600 53.100 129.000 53.200 ;
        RECT 122.200 52.800 123.400 53.100 ;
        RECT 126.200 52.800 129.000 53.100 ;
        RECT 137.400 53.100 137.800 53.200 ;
        RECT 138.200 53.100 138.600 53.200 ;
        RECT 137.400 52.800 138.600 53.100 ;
        RECT 87.000 52.200 87.300 52.800 ;
        RECT 126.200 52.200 126.500 52.800 ;
        RECT 11.800 52.100 12.200 52.200 ;
        RECT 18.200 52.100 18.600 52.200 ;
        RECT 20.600 52.100 21.000 52.200 ;
        RECT 11.800 51.800 21.000 52.100 ;
        RECT 43.800 52.100 44.200 52.200 ;
        RECT 46.200 52.100 46.600 52.200 ;
        RECT 43.800 51.800 46.600 52.100 ;
        RECT 63.800 52.100 64.200 52.200 ;
        RECT 72.600 52.100 73.000 52.200 ;
        RECT 63.800 51.800 73.000 52.100 ;
        RECT 78.200 52.100 78.600 52.200 ;
        RECT 83.800 52.100 84.200 52.200 ;
        RECT 85.400 52.100 85.800 52.200 ;
        RECT 78.200 51.800 85.800 52.100 ;
        RECT 87.000 51.800 87.400 52.200 ;
        RECT 90.200 52.100 90.600 52.200 ;
        RECT 95.800 52.100 96.200 52.200 ;
        RECT 104.600 52.100 105.000 52.200 ;
        RECT 89.400 51.800 96.200 52.100 ;
        RECT 96.600 51.800 105.000 52.100 ;
        RECT 105.400 52.100 105.800 52.200 ;
        RECT 119.800 52.100 120.200 52.200 ;
        RECT 105.400 51.800 120.200 52.100 ;
        RECT 126.200 51.800 126.600 52.200 ;
        RECT 131.000 52.100 131.400 52.200 ;
        RECT 132.600 52.100 133.000 52.200 ;
        RECT 131.000 51.800 133.000 52.100 ;
        RECT 96.600 51.200 96.900 51.800 ;
        RECT 58.200 51.100 58.600 51.200 ;
        RECT 82.200 51.100 82.600 51.200 ;
        RECT 58.200 50.800 82.600 51.100 ;
        RECT 87.000 51.100 87.400 51.200 ;
        RECT 91.800 51.100 92.200 51.200 ;
        RECT 87.000 50.800 92.200 51.100 ;
        RECT 92.600 51.100 93.000 51.200 ;
        RECT 93.400 51.100 93.800 51.200 ;
        RECT 92.600 50.800 93.800 51.100 ;
        RECT 96.600 50.800 97.000 51.200 ;
        RECT 111.000 51.100 111.400 51.200 ;
        RECT 127.000 51.100 127.400 51.200 ;
        RECT 133.400 51.100 133.800 51.200 ;
        RECT 111.000 50.800 133.800 51.100 ;
        RECT 63.000 50.100 63.400 50.200 ;
        RECT 69.400 50.100 69.800 50.200 ;
        RECT 63.000 49.800 69.800 50.100 ;
        RECT 83.000 50.100 83.400 50.200 ;
        RECT 98.200 50.100 98.600 50.200 ;
        RECT 83.000 49.800 98.600 50.100 ;
        RECT 103.000 50.100 103.400 50.200 ;
        RECT 111.800 50.100 112.200 50.200 ;
        RECT 103.000 49.800 112.200 50.100 ;
        RECT 43.000 48.800 43.400 49.200 ;
        RECT 44.600 48.800 45.000 49.200 ;
        RECT 59.000 49.100 59.400 49.200 ;
        RECT 80.600 49.100 81.000 49.200 ;
        RECT 97.400 49.100 97.800 49.200 ;
        RECT 59.000 48.800 81.000 49.100 ;
        RECT 81.400 48.800 97.800 49.100 ;
        RECT 98.200 49.100 98.600 49.200 ;
        RECT 103.000 49.100 103.400 49.200 ;
        RECT 107.800 49.100 108.200 49.200 ;
        RECT 98.200 48.800 108.200 49.100 ;
        RECT 115.000 49.100 115.400 49.200 ;
        RECT 123.800 49.100 124.200 49.200 ;
        RECT 131.800 49.100 132.200 49.200 ;
        RECT 135.000 49.100 135.400 49.200 ;
        RECT 115.000 48.800 135.400 49.100 ;
        RECT 137.400 48.800 137.800 49.200 ;
        RECT 145.400 49.100 145.800 49.200 ;
        RECT 147.000 49.100 147.400 49.200 ;
        RECT 145.400 48.800 147.400 49.100 ;
        RECT 16.600 47.800 17.000 48.200 ;
        RECT 35.000 48.100 35.400 48.200 ;
        RECT 38.200 48.100 38.600 48.200 ;
        RECT 35.000 47.800 38.600 48.100 ;
        RECT 39.800 48.100 40.200 48.200 ;
        RECT 43.000 48.100 43.300 48.800 ;
        RECT 39.800 47.800 43.300 48.100 ;
        RECT 44.600 48.200 44.900 48.800 ;
        RECT 81.400 48.200 81.700 48.800 ;
        RECT 137.400 48.200 137.700 48.800 ;
        RECT 44.600 47.800 45.000 48.200 ;
        RECT 56.600 47.800 57.000 48.200 ;
        RECT 60.600 48.100 61.000 48.200 ;
        RECT 73.400 48.100 73.800 48.200 ;
        RECT 60.600 47.800 73.800 48.100 ;
        RECT 81.400 47.800 81.800 48.200 ;
        RECT 84.600 47.800 85.000 48.200 ;
        RECT 86.200 48.100 86.600 48.200 ;
        RECT 87.000 48.100 87.400 48.200 ;
        RECT 86.200 47.800 87.400 48.100 ;
        RECT 88.600 48.100 89.000 48.200 ;
        RECT 94.200 48.100 94.600 48.200 ;
        RECT 98.200 48.100 98.600 48.200 ;
        RECT 88.600 47.800 98.600 48.100 ;
        RECT 99.000 48.100 99.400 48.200 ;
        RECT 111.000 48.100 111.400 48.200 ;
        RECT 115.000 48.100 115.400 48.200 ;
        RECT 99.000 47.800 115.400 48.100 ;
        RECT 137.400 47.800 137.800 48.200 ;
        RECT 11.000 47.100 11.400 47.200 ;
        RECT 16.600 47.100 16.900 47.800 ;
        RECT 11.000 46.800 16.900 47.100 ;
        RECT 23.000 46.800 23.400 47.200 ;
        RECT 42.200 47.100 42.600 47.200 ;
        RECT 47.800 47.100 48.200 47.200 ;
        RECT 56.600 47.100 56.900 47.800 ;
        RECT 42.200 46.800 56.900 47.100 ;
        RECT 66.200 47.100 66.600 47.200 ;
        RECT 84.600 47.100 84.900 47.800 ;
        RECT 66.200 46.800 84.900 47.100 ;
        RECT 86.200 47.100 86.600 47.200 ;
        RECT 90.200 47.100 90.600 47.200 ;
        RECT 86.200 46.800 90.600 47.100 ;
        RECT 97.400 47.100 97.800 47.200 ;
        RECT 100.600 47.100 101.000 47.200 ;
        RECT 107.000 47.100 107.400 47.200 ;
        RECT 97.400 46.800 107.400 47.100 ;
        RECT 115.000 46.800 115.400 47.200 ;
        RECT 116.600 47.100 117.000 47.200 ;
        RECT 117.400 47.100 117.800 47.200 ;
        RECT 120.600 47.100 121.000 47.200 ;
        RECT 116.600 46.800 121.000 47.100 ;
        RECT 125.400 47.100 125.800 47.200 ;
        RECT 131.000 47.100 131.400 47.200 ;
        RECT 125.400 46.800 131.400 47.100 ;
        RECT 138.200 47.100 138.600 47.200 ;
        RECT 139.800 47.100 140.200 47.200 ;
        RECT 145.400 47.100 145.800 47.200 ;
        RECT 148.600 47.100 149.000 47.200 ;
        RECT 138.200 46.800 149.000 47.100 ;
        RECT 6.200 46.100 6.600 46.200 ;
        RECT 9.400 46.100 9.800 46.200 ;
        RECT 6.200 45.800 9.800 46.100 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 23.000 46.100 23.300 46.800 ;
        RECT 27.800 46.100 28.200 46.200 ;
        RECT 14.200 45.800 20.100 46.100 ;
        RECT 23.000 45.800 28.200 46.100 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 35.000 46.100 35.400 46.200 ;
        RECT 38.200 46.100 38.600 46.200 ;
        RECT 31.800 45.800 38.600 46.100 ;
        RECT 39.000 46.100 39.400 46.200 ;
        RECT 45.400 46.100 45.800 46.200 ;
        RECT 39.000 45.800 45.800 46.100 ;
        RECT 47.000 46.100 47.400 46.200 ;
        RECT 48.600 46.100 49.000 46.200 ;
        RECT 47.000 45.800 49.000 46.100 ;
        RECT 61.400 46.100 61.800 46.200 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 67.800 46.100 68.200 46.200 ;
        RECT 61.400 45.800 68.200 46.100 ;
        RECT 69.400 46.100 69.800 46.200 ;
        RECT 75.000 46.100 75.400 46.200 ;
        RECT 69.400 45.800 75.400 46.100 ;
        RECT 77.400 46.100 77.800 46.200 ;
        RECT 87.800 46.100 88.200 46.200 ;
        RECT 77.400 45.800 88.200 46.100 ;
        RECT 89.400 46.100 89.800 46.200 ;
        RECT 96.600 46.100 97.000 46.200 ;
        RECT 89.400 45.800 97.000 46.100 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 110.200 46.100 110.600 46.200 ;
        RECT 98.200 45.800 110.600 46.100 ;
        RECT 115.000 46.100 115.300 46.800 ;
        RECT 117.400 46.100 117.800 46.200 ;
        RECT 119.000 46.100 119.400 46.200 ;
        RECT 115.000 45.800 119.400 46.100 ;
        RECT 136.600 46.100 137.000 46.200 ;
        RECT 137.400 46.100 137.800 46.200 ;
        RECT 141.400 46.100 141.800 46.200 ;
        RECT 147.000 46.100 147.400 46.200 ;
        RECT 136.600 45.800 147.400 46.100 ;
        RECT 19.800 45.200 20.100 45.800 ;
        RECT 3.000 45.100 3.400 45.200 ;
        RECT 7.800 45.100 8.200 45.200 ;
        RECT 3.000 44.800 8.200 45.100 ;
        RECT 19.800 44.800 20.200 45.200 ;
        RECT 38.200 45.100 38.600 45.200 ;
        RECT 40.600 45.100 41.000 45.200 ;
        RECT 38.200 44.800 41.000 45.100 ;
        RECT 43.000 45.100 43.400 45.200 ;
        RECT 46.200 45.100 46.600 45.200 ;
        RECT 79.000 45.100 79.400 45.200 ;
        RECT 80.600 45.100 81.000 45.200 ;
        RECT 43.000 44.800 46.600 45.100 ;
        RECT 78.200 44.800 81.000 45.100 ;
        RECT 82.200 45.100 82.600 45.200 ;
        RECT 85.400 45.100 85.800 45.200 ;
        RECT 91.000 45.100 91.400 45.200 ;
        RECT 93.400 45.100 93.800 45.200 ;
        RECT 82.200 44.800 93.800 45.100 ;
        RECT 95.800 45.100 96.200 45.200 ;
        RECT 103.800 45.100 104.200 45.200 ;
        RECT 105.400 45.100 105.800 45.200 ;
        RECT 95.800 44.800 105.800 45.100 ;
        RECT 139.800 45.100 140.200 45.200 ;
        RECT 143.000 45.100 143.400 45.200 ;
        RECT 139.800 44.800 143.400 45.100 ;
        RECT 144.600 44.800 145.000 45.200 ;
        RECT 144.600 44.200 144.900 44.800 ;
        RECT 75.000 44.100 75.400 44.200 ;
        RECT 122.200 44.100 122.600 44.200 ;
        RECT 126.200 44.100 126.600 44.200 ;
        RECT 132.600 44.100 133.000 44.200 ;
        RECT 135.800 44.100 136.200 44.200 ;
        RECT 75.000 43.800 136.200 44.100 ;
        RECT 144.600 44.100 145.000 44.200 ;
        RECT 147.000 44.100 147.400 44.200 ;
        RECT 144.600 43.800 147.400 44.100 ;
        RECT 52.600 43.100 53.000 43.200 ;
        RECT 59.800 43.100 60.200 43.200 ;
        RECT 52.600 42.800 60.200 43.100 ;
        RECT 64.600 43.100 65.000 43.200 ;
        RECT 83.800 43.100 84.200 43.200 ;
        RECT 87.800 43.100 88.200 43.200 ;
        RECT 64.600 42.800 88.200 43.100 ;
        RECT 17.400 42.100 17.800 42.200 ;
        RECT 18.200 42.100 18.600 42.200 ;
        RECT 17.400 41.800 18.600 42.100 ;
        RECT 79.800 42.100 80.200 42.200 ;
        RECT 86.200 42.100 86.600 42.200 ;
        RECT 79.800 41.800 86.600 42.100 ;
        RECT 135.800 42.100 136.200 42.200 ;
        RECT 137.400 42.100 137.800 42.200 ;
        RECT 138.200 42.100 138.600 42.200 ;
        RECT 135.800 41.800 138.600 42.100 ;
        RECT 63.800 41.100 64.200 41.200 ;
        RECT 65.400 41.100 65.800 41.200 ;
        RECT 63.800 40.800 65.800 41.100 ;
        RECT 20.600 39.100 21.000 39.200 ;
        RECT 22.200 39.100 22.600 39.200 ;
        RECT 20.600 38.800 22.600 39.100 ;
        RECT 27.000 39.100 27.400 39.200 ;
        RECT 27.800 39.100 28.200 39.200 ;
        RECT 27.000 38.800 28.200 39.100 ;
        RECT 80.600 38.100 81.000 38.200 ;
        RECT 81.400 38.100 81.800 38.200 ;
        RECT 83.800 38.100 84.200 38.200 ;
        RECT 80.600 37.800 84.200 38.100 ;
        RECT 7.000 36.800 7.400 37.200 ;
        RECT 45.400 36.800 45.800 37.200 ;
        RECT 87.800 37.100 88.200 37.200 ;
        RECT 113.400 37.100 113.800 37.200 ;
        RECT 87.800 36.800 113.800 37.100 ;
        RECT 146.200 36.800 146.600 37.200 ;
        RECT 7.000 36.100 7.300 36.800 ;
        RECT 9.400 36.100 9.800 36.200 ;
        RECT 7.000 35.800 9.800 36.100 ;
        RECT 15.800 36.100 16.200 36.200 ;
        RECT 21.400 36.100 21.800 36.200 ;
        RECT 15.800 35.800 21.800 36.100 ;
        RECT 37.400 35.800 37.800 36.200 ;
        RECT 42.200 36.100 42.600 36.200 ;
        RECT 45.400 36.100 45.700 36.800 ;
        RECT 146.200 36.200 146.500 36.800 ;
        RECT 48.600 36.100 49.000 36.200 ;
        RECT 42.200 35.800 49.000 36.100 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 75.000 36.100 75.400 36.200 ;
        RECT 76.600 36.100 77.000 36.200 ;
        RECT 80.600 36.100 81.000 36.200 ;
        RECT 75.000 35.800 81.000 36.100 ;
        RECT 85.400 36.100 85.800 36.200 ;
        RECT 88.600 36.100 89.000 36.200 ;
        RECT 85.400 35.800 89.000 36.100 ;
        RECT 91.000 36.100 91.400 36.200 ;
        RECT 97.400 36.100 97.800 36.200 ;
        RECT 91.000 35.800 97.800 36.100 ;
        RECT 112.600 36.100 113.000 36.200 ;
        RECT 118.200 36.100 118.600 36.200 ;
        RECT 112.600 35.800 118.600 36.100 ;
        RECT 124.600 36.100 125.000 36.200 ;
        RECT 131.000 36.100 131.400 36.200 ;
        RECT 124.600 35.800 131.400 36.100 ;
        RECT 133.400 35.800 133.800 36.200 ;
        RECT 136.600 36.100 137.000 36.200 ;
        RECT 139.000 36.100 139.400 36.200 ;
        RECT 136.600 35.800 139.400 36.100 ;
        RECT 146.200 35.800 146.600 36.200 ;
        RECT 3.000 35.100 3.400 35.200 ;
        RECT 11.000 35.100 11.400 35.200 ;
        RECT 3.000 34.800 11.400 35.100 ;
        RECT 12.600 35.100 13.000 35.200 ;
        RECT 18.200 35.100 18.600 35.200 ;
        RECT 12.600 34.800 18.600 35.100 ;
        RECT 37.400 35.100 37.700 35.800 ;
        RECT 67.000 35.100 67.300 35.800 ;
        RECT 37.400 34.800 67.300 35.100 ;
        RECT 80.600 35.100 81.000 35.200 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 86.200 35.100 86.600 35.200 ;
        RECT 80.600 34.800 86.600 35.100 ;
        RECT 92.600 35.100 93.000 35.200 ;
        RECT 105.400 35.100 105.800 35.200 ;
        RECT 109.400 35.100 109.800 35.200 ;
        RECT 92.600 34.800 93.700 35.100 ;
        RECT 105.400 34.800 109.800 35.100 ;
        RECT 111.800 35.100 112.200 35.200 ;
        RECT 115.000 35.100 115.400 35.200 ;
        RECT 111.800 34.800 115.400 35.100 ;
        RECT 123.000 35.100 123.400 35.200 ;
        RECT 126.200 35.100 126.600 35.200 ;
        RECT 127.800 35.100 128.200 35.200 ;
        RECT 123.000 34.800 128.200 35.100 ;
        RECT 133.400 35.100 133.700 35.800 ;
        RECT 138.200 35.100 138.600 35.200 ;
        RECT 133.400 34.800 138.600 35.100 ;
        RECT 143.000 35.100 143.400 35.200 ;
        RECT 143.800 35.100 144.200 35.200 ;
        RECT 143.000 34.800 144.200 35.100 ;
        RECT 93.400 34.200 93.700 34.800 ;
        RECT 47.000 34.100 47.400 34.200 ;
        RECT 60.600 34.100 61.000 34.200 ;
        RECT 72.600 34.100 73.000 34.200 ;
        RECT 73.400 34.100 73.800 34.200 ;
        RECT 47.000 33.800 54.500 34.100 ;
        RECT 60.600 33.800 65.700 34.100 ;
        RECT 72.600 33.800 73.800 34.100 ;
        RECT 76.600 34.100 77.000 34.200 ;
        RECT 87.800 34.100 88.200 34.200 ;
        RECT 76.600 33.800 88.200 34.100 ;
        RECT 89.400 34.100 89.800 34.200 ;
        RECT 91.800 34.100 92.200 34.200 ;
        RECT 89.400 33.800 92.200 34.100 ;
        RECT 93.400 33.800 93.800 34.200 ;
        RECT 103.000 34.100 103.400 34.200 ;
        RECT 107.000 34.100 107.400 34.200 ;
        RECT 111.000 34.100 111.400 34.200 ;
        RECT 103.000 33.800 111.400 34.100 ;
        RECT 123.800 34.100 124.200 34.200 ;
        RECT 125.400 34.100 125.800 34.200 ;
        RECT 123.800 33.800 125.800 34.100 ;
        RECT 139.000 34.100 139.400 34.200 ;
        RECT 140.600 34.100 141.000 34.200 ;
        RECT 139.000 33.800 141.000 34.100 ;
        RECT 54.200 33.200 54.500 33.800 ;
        RECT 65.400 33.200 65.700 33.800 ;
        RECT 54.200 32.800 54.600 33.200 ;
        RECT 65.400 32.800 65.800 33.200 ;
        RECT 77.400 33.100 77.800 33.200 ;
        RECT 82.200 33.100 82.600 33.200 ;
        RECT 77.400 32.800 82.600 33.100 ;
        RECT 83.000 33.100 83.400 33.200 ;
        RECT 87.000 33.100 87.400 33.200 ;
        RECT 91.000 33.100 91.400 33.200 ;
        RECT 97.400 33.100 97.800 33.200 ;
        RECT 112.600 33.100 113.000 33.200 ;
        RECT 83.000 32.800 89.700 33.100 ;
        RECT 91.000 32.800 97.800 33.100 ;
        RECT 107.000 32.800 113.000 33.100 ;
        RECT 125.400 32.800 125.800 33.200 ;
        RECT 134.200 33.100 134.600 33.200 ;
        RECT 142.200 33.100 142.600 33.200 ;
        RECT 134.200 32.800 142.600 33.100 ;
        RECT 89.400 32.200 89.700 32.800 ;
        RECT 107.000 32.200 107.300 32.800 ;
        RECT 125.400 32.200 125.700 32.800 ;
        RECT 74.200 32.100 74.600 32.200 ;
        RECT 79.000 32.100 79.400 32.200 ;
        RECT 74.200 31.800 79.400 32.100 ;
        RECT 89.400 31.800 89.800 32.200 ;
        RECT 93.400 32.100 93.800 32.200 ;
        RECT 107.000 32.100 107.400 32.200 ;
        RECT 93.400 31.800 107.400 32.100 ;
        RECT 125.400 32.100 125.800 32.200 ;
        RECT 141.400 32.100 141.800 32.200 ;
        RECT 125.400 31.800 141.800 32.100 ;
        RECT 71.000 31.100 71.400 31.200 ;
        RECT 90.200 31.100 90.600 31.200 ;
        RECT 95.800 31.100 96.200 31.200 ;
        RECT 71.000 30.800 96.200 31.100 ;
        RECT 110.200 31.100 110.600 31.200 ;
        RECT 113.400 31.100 113.800 31.200 ;
        RECT 110.200 30.800 113.800 31.100 ;
        RECT 144.600 31.100 145.000 31.200 ;
        RECT 147.000 31.100 147.400 31.200 ;
        RECT 144.600 30.800 147.400 31.100 ;
        RECT 84.600 30.100 85.000 30.200 ;
        RECT 86.200 30.100 86.600 30.200 ;
        RECT 114.200 30.100 114.600 30.200 ;
        RECT 84.600 29.800 86.600 30.100 ;
        RECT 111.000 29.800 114.600 30.100 ;
        RECT 147.000 30.100 147.400 30.200 ;
        RECT 151.000 30.100 151.400 30.200 ;
        RECT 147.000 29.800 151.400 30.100 ;
        RECT 111.000 29.200 111.300 29.800 ;
        RECT 39.800 29.100 40.200 29.200 ;
        RECT 40.600 29.100 41.000 29.200 ;
        RECT 39.800 28.800 41.000 29.100 ;
        RECT 51.000 29.100 51.400 29.200 ;
        RECT 51.800 29.100 52.200 29.200 ;
        RECT 51.000 28.800 52.200 29.100 ;
        RECT 63.000 29.100 63.400 29.200 ;
        RECT 71.800 29.100 72.200 29.200 ;
        RECT 89.400 29.100 89.800 29.200 ;
        RECT 90.200 29.100 90.600 29.200 ;
        RECT 63.000 28.800 90.600 29.100 ;
        RECT 103.000 29.100 103.400 29.200 ;
        RECT 111.000 29.100 111.400 29.200 ;
        RECT 103.000 28.800 111.400 29.100 ;
        RECT 115.000 29.100 115.400 29.200 ;
        RECT 116.600 29.100 117.000 29.200 ;
        RECT 115.000 28.800 117.000 29.100 ;
        RECT 129.400 29.100 129.800 29.200 ;
        RECT 131.000 29.100 131.400 29.200 ;
        RECT 129.400 28.800 131.400 29.100 ;
        RECT 33.400 27.800 33.800 28.200 ;
        RECT 51.000 28.100 51.400 28.200 ;
        RECT 58.200 28.100 58.600 28.200 ;
        RECT 51.000 27.800 58.600 28.100 ;
        RECT 77.400 27.800 77.800 28.200 ;
        RECT 94.200 28.100 94.600 28.200 ;
        RECT 100.600 28.100 101.000 28.200 ;
        RECT 104.600 28.100 105.000 28.200 ;
        RECT 85.400 27.800 105.000 28.100 ;
        RECT 112.600 28.100 113.000 28.200 ;
        RECT 119.000 28.100 119.400 28.200 ;
        RECT 112.600 27.800 119.400 28.100 ;
        RECT 121.400 28.100 121.800 28.200 ;
        RECT 125.400 28.100 125.800 28.200 ;
        RECT 121.400 27.800 125.800 28.100 ;
        RECT 127.000 28.100 127.400 28.200 ;
        RECT 133.400 28.100 133.800 28.200 ;
        RECT 127.000 27.800 133.800 28.100 ;
        RECT 3.800 27.100 4.200 27.200 ;
        RECT 7.000 27.100 7.400 27.200 ;
        RECT 3.800 26.800 7.400 27.100 ;
        RECT 20.600 27.100 21.000 27.200 ;
        RECT 21.400 27.100 21.800 27.200 ;
        RECT 31.000 27.100 31.400 27.200 ;
        RECT 33.400 27.100 33.700 27.800 ;
        RECT 20.600 26.800 33.700 27.100 ;
        RECT 47.800 26.800 48.200 27.200 ;
        RECT 77.400 27.100 77.700 27.800 ;
        RECT 85.400 27.200 85.700 27.800 ;
        RECT 83.000 27.100 83.400 27.200 ;
        RECT 77.400 26.800 83.400 27.100 ;
        RECT 85.400 26.800 85.800 27.200 ;
        RECT 87.000 26.800 87.400 27.200 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 103.000 27.100 103.400 27.200 ;
        RECT 95.000 26.800 103.400 27.100 ;
        RECT 107.800 27.100 108.200 27.200 ;
        RECT 111.800 27.100 112.200 27.200 ;
        RECT 107.800 26.800 112.200 27.100 ;
        RECT 117.400 27.100 117.800 27.200 ;
        RECT 119.800 27.100 120.200 27.200 ;
        RECT 125.400 27.100 125.800 27.200 ;
        RECT 128.600 27.100 129.000 27.200 ;
        RECT 117.400 26.800 129.000 27.100 ;
        RECT 131.000 27.100 131.400 27.200 ;
        RECT 131.800 27.100 132.200 27.200 ;
        RECT 136.600 27.100 137.000 27.200 ;
        RECT 131.000 26.800 137.000 27.100 ;
        RECT 143.800 27.100 144.200 27.200 ;
        RECT 145.400 27.100 145.800 27.200 ;
        RECT 143.800 26.800 145.800 27.100 ;
        RECT 148.600 26.800 149.000 27.200 ;
        RECT 23.800 26.200 24.100 26.800 ;
        RECT 9.400 25.800 16.100 26.100 ;
        RECT 23.800 25.800 24.200 26.200 ;
        RECT 30.200 26.100 30.600 26.200 ;
        RECT 47.800 26.100 48.100 26.800 ;
        RECT 57.400 26.100 57.800 26.200 ;
        RECT 30.200 25.800 35.300 26.100 ;
        RECT 47.800 25.800 57.800 26.100 ;
        RECT 83.800 26.100 84.200 26.200 ;
        RECT 87.000 26.100 87.300 26.800 ;
        RECT 83.800 25.800 87.300 26.100 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 99.000 26.100 99.400 26.200 ;
        RECT 97.400 25.800 99.400 26.100 ;
        RECT 106.200 26.100 106.600 26.200 ;
        RECT 109.400 26.100 109.800 26.200 ;
        RECT 106.200 25.800 109.800 26.100 ;
        RECT 110.200 26.100 110.600 26.200 ;
        RECT 129.400 26.100 129.800 26.200 ;
        RECT 110.200 25.800 129.800 26.100 ;
        RECT 131.000 26.100 131.400 26.200 ;
        RECT 133.400 26.100 133.800 26.200 ;
        RECT 138.200 26.100 138.600 26.200 ;
        RECT 131.000 25.800 138.600 26.100 ;
        RECT 143.800 26.100 144.200 26.200 ;
        RECT 148.600 26.100 148.900 26.800 ;
        RECT 143.800 25.800 148.900 26.100 ;
        RECT 9.400 25.200 9.700 25.800 ;
        RECT 15.800 25.200 16.100 25.800 ;
        RECT 35.000 25.200 35.300 25.800 ;
        RECT 9.400 24.800 9.800 25.200 ;
        RECT 15.800 24.800 16.200 25.200 ;
        RECT 35.000 24.800 35.400 25.200 ;
        RECT 87.800 25.100 88.200 25.200 ;
        RECT 91.000 25.100 91.400 25.200 ;
        RECT 87.800 24.800 91.400 25.100 ;
        RECT 99.800 25.100 100.200 25.200 ;
        RECT 104.600 25.100 105.000 25.200 ;
        RECT 107.000 25.100 107.400 25.200 ;
        RECT 99.800 24.800 107.400 25.100 ;
        RECT 131.800 25.100 132.200 25.200 ;
        RECT 137.400 25.100 137.800 25.200 ;
        RECT 131.800 24.800 137.800 25.100 ;
        RECT 139.800 25.100 140.200 25.200 ;
        RECT 143.000 25.100 143.400 25.200 ;
        RECT 139.800 24.800 143.400 25.100 ;
        RECT 145.400 25.100 145.800 25.200 ;
        RECT 146.200 25.100 146.600 25.200 ;
        RECT 145.400 24.800 146.600 25.100 ;
        RECT 6.200 24.100 6.600 24.200 ;
        RECT 14.200 24.100 14.600 24.200 ;
        RECT 6.200 23.800 14.600 24.100 ;
        RECT 26.200 24.100 26.600 24.200 ;
        RECT 55.800 24.100 56.200 24.200 ;
        RECT 26.200 23.800 56.200 24.100 ;
        RECT 119.000 24.100 119.400 24.200 ;
        RECT 135.000 24.100 135.400 24.200 ;
        RECT 119.000 23.800 135.400 24.100 ;
        RECT 141.400 24.100 141.800 24.200 ;
        RECT 144.600 24.100 145.000 24.200 ;
        RECT 141.400 23.800 145.000 24.100 ;
        RECT 8.600 23.100 9.000 23.200 ;
        RECT 15.800 23.100 16.200 23.200 ;
        RECT 8.600 22.800 16.200 23.100 ;
        RECT 136.600 23.100 137.000 23.200 ;
        RECT 140.600 23.100 141.000 23.200 ;
        RECT 136.600 22.800 141.000 23.100 ;
        RECT 9.400 22.100 9.800 22.200 ;
        RECT 44.600 22.100 45.000 22.200 ;
        RECT 9.400 21.800 45.000 22.100 ;
        RECT 128.600 22.100 129.000 22.200 ;
        RECT 139.000 22.100 139.400 22.200 ;
        RECT 128.600 21.800 139.400 22.100 ;
        RECT 105.400 20.100 105.800 20.200 ;
        RECT 115.800 20.100 116.200 20.200 ;
        RECT 105.400 19.800 116.200 20.100 ;
        RECT 69.400 19.100 69.800 19.200 ;
        RECT 82.200 19.100 82.600 19.200 ;
        RECT 111.000 19.100 111.400 19.200 ;
        RECT 124.600 19.100 125.000 19.200 ;
        RECT 69.400 18.800 82.600 19.100 ;
        RECT 104.600 18.800 125.000 19.100 ;
        RECT 146.200 19.100 146.600 19.200 ;
        RECT 146.200 18.800 148.100 19.100 ;
        RECT 104.600 18.200 104.900 18.800 ;
        RECT 147.800 18.200 148.100 18.800 ;
        RECT 70.200 18.100 70.600 18.200 ;
        RECT 76.600 18.100 77.000 18.200 ;
        RECT 70.200 17.800 77.000 18.100 ;
        RECT 104.600 17.800 105.000 18.200 ;
        RECT 109.400 17.800 109.800 18.200 ;
        RECT 147.800 17.800 148.200 18.200 ;
        RECT 42.200 16.800 42.600 17.200 ;
        RECT 61.400 17.100 61.800 17.200 ;
        RECT 61.400 16.800 72.900 17.100 ;
        RECT 42.200 16.100 42.500 16.800 ;
        RECT 72.600 16.200 72.900 16.800 ;
        RECT 76.600 16.800 77.000 17.200 ;
        RECT 92.600 17.100 93.000 17.200 ;
        RECT 95.000 17.100 95.400 17.200 ;
        RECT 92.600 16.800 95.400 17.100 ;
        RECT 102.200 17.100 102.600 17.200 ;
        RECT 103.000 17.100 103.400 17.200 ;
        RECT 102.200 16.800 103.400 17.100 ;
        RECT 109.400 17.100 109.700 17.800 ;
        RECT 111.800 17.100 112.200 17.200 ;
        RECT 109.400 16.800 112.200 17.100 ;
        RECT 122.200 17.100 122.600 17.200 ;
        RECT 126.200 17.100 126.600 17.200 ;
        RECT 122.200 16.800 126.600 17.100 ;
        RECT 148.600 16.800 149.000 17.200 ;
        RECT 47.000 16.100 47.400 16.200 ;
        RECT 49.400 16.100 49.800 16.200 ;
        RECT 42.200 15.800 49.800 16.100 ;
        RECT 72.600 15.800 73.000 16.200 ;
        RECT 76.600 16.100 76.900 16.800 ;
        RECT 148.600 16.200 148.900 16.800 ;
        RECT 85.400 16.100 85.800 16.200 ;
        RECT 76.600 15.800 85.800 16.100 ;
        RECT 93.400 16.100 93.800 16.200 ;
        RECT 95.000 16.100 95.400 16.200 ;
        RECT 106.200 16.100 106.600 16.200 ;
        RECT 93.400 15.800 106.600 16.100 ;
        RECT 107.000 16.100 107.400 16.200 ;
        RECT 109.400 16.100 109.800 16.200 ;
        RECT 115.000 16.100 115.400 16.200 ;
        RECT 107.000 15.800 115.400 16.100 ;
        RECT 125.400 16.100 125.800 16.200 ;
        RECT 126.200 16.100 126.600 16.200 ;
        RECT 125.400 15.800 126.600 16.100 ;
        RECT 137.400 15.800 137.800 16.200 ;
        RECT 148.600 15.800 149.000 16.200 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 44.600 15.100 45.000 15.200 ;
        RECT 41.400 14.800 45.000 15.100 ;
        RECT 48.600 15.100 49.000 15.200 ;
        RECT 60.600 15.100 61.000 15.200 ;
        RECT 73.400 15.100 73.800 15.200 ;
        RECT 77.400 15.100 77.800 15.200 ;
        RECT 48.600 14.800 54.500 15.100 ;
        RECT 60.600 14.800 64.900 15.100 ;
        RECT 73.400 14.800 77.800 15.100 ;
        RECT 83.800 15.100 84.200 15.200 ;
        RECT 84.600 15.100 85.000 15.200 ;
        RECT 94.200 15.100 94.600 15.200 ;
        RECT 83.800 14.800 85.000 15.100 ;
        RECT 90.200 14.800 94.600 15.100 ;
        RECT 105.400 15.100 105.800 15.200 ;
        RECT 110.200 15.100 110.600 15.200 ;
        RECT 115.800 15.100 116.200 15.200 ;
        RECT 105.400 14.800 106.500 15.100 ;
        RECT 110.200 14.800 116.200 15.100 ;
        RECT 123.800 15.100 124.200 15.200 ;
        RECT 127.000 15.100 127.400 15.200 ;
        RECT 123.800 14.800 127.400 15.100 ;
        RECT 132.600 15.100 133.000 15.200 ;
        RECT 137.400 15.100 137.700 15.800 ;
        RECT 132.600 14.800 137.700 15.100 ;
        RECT 43.800 14.200 44.100 14.800 ;
        RECT 54.200 14.200 54.500 14.800 ;
        RECT 64.600 14.200 64.900 14.800 ;
        RECT 90.200 14.200 90.500 14.800 ;
        RECT 43.800 13.800 44.200 14.200 ;
        RECT 54.200 13.800 54.600 14.200 ;
        RECT 57.400 14.100 57.800 14.200 ;
        RECT 63.800 14.100 64.200 14.200 ;
        RECT 57.400 13.800 64.200 14.100 ;
        RECT 64.600 13.800 65.000 14.200 ;
        RECT 75.000 14.100 75.400 14.200 ;
        RECT 76.600 14.100 77.000 14.200 ;
        RECT 75.000 13.800 77.000 14.100 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 90.200 14.100 90.600 14.200 ;
        RECT 82.200 13.800 90.600 14.100 ;
        RECT 91.800 13.800 92.200 14.200 ;
        RECT 97.400 14.100 97.800 14.200 ;
        RECT 102.200 14.100 102.600 14.200 ;
        RECT 107.800 14.100 108.200 14.200 ;
        RECT 114.200 14.100 114.600 14.200 ;
        RECT 97.400 13.800 114.600 14.100 ;
        RECT 120.600 14.100 121.000 14.200 ;
        RECT 126.200 14.100 126.600 14.200 ;
        RECT 120.600 13.800 126.600 14.100 ;
        RECT 147.800 14.100 148.200 14.200 ;
        RECT 150.200 14.100 150.600 14.200 ;
        RECT 147.800 13.800 150.600 14.100 ;
        RECT 45.400 13.100 45.800 13.200 ;
        RECT 46.200 13.100 46.600 13.200 ;
        RECT 47.800 13.100 48.200 13.200 ;
        RECT 45.400 12.800 48.200 13.100 ;
        RECT 79.800 12.800 80.200 13.200 ;
        RECT 83.000 13.100 83.400 13.200 ;
        RECT 85.400 13.100 85.800 13.200 ;
        RECT 83.000 12.800 85.800 13.100 ;
        RECT 91.800 13.100 92.100 13.800 ;
        RECT 96.600 13.100 97.000 13.200 ;
        RECT 123.000 13.100 123.400 13.200 ;
        RECT 91.800 12.800 97.000 13.100 ;
        RECT 121.400 12.800 123.400 13.100 ;
        RECT 145.400 13.100 145.800 13.200 ;
        RECT 147.000 13.100 147.400 13.200 ;
        RECT 145.400 12.800 147.400 13.100 ;
        RECT 11.800 12.100 12.200 12.200 ;
        RECT 14.200 12.100 14.600 12.200 ;
        RECT 11.800 11.800 14.600 12.100 ;
        RECT 15.000 12.100 15.400 12.200 ;
        RECT 25.400 12.100 25.800 12.200 ;
        RECT 15.000 11.800 25.800 12.100 ;
        RECT 79.800 12.100 80.100 12.800 ;
        RECT 121.400 12.200 121.700 12.800 ;
        RECT 87.800 12.100 88.200 12.200 ;
        RECT 79.800 11.800 88.200 12.100 ;
        RECT 121.400 11.800 121.800 12.200 ;
        RECT 24.600 9.100 25.000 9.200 ;
        RECT 27.000 9.100 27.400 9.200 ;
        RECT 24.600 8.800 27.400 9.100 ;
        RECT 44.600 8.100 45.000 8.200 ;
        RECT 54.200 8.100 54.600 8.200 ;
        RECT 44.600 7.800 54.600 8.100 ;
        RECT 71.800 7.800 72.200 8.200 ;
        RECT 99.800 8.100 100.200 8.200 ;
        RECT 111.800 8.100 112.200 8.200 ;
        RECT 123.800 8.100 124.200 8.200 ;
        RECT 135.800 8.100 136.200 8.200 ;
        RECT 99.800 7.800 136.200 8.100 ;
        RECT 7.000 7.100 7.400 7.200 ;
        RECT 11.800 7.100 12.200 7.200 ;
        RECT 7.000 6.800 12.200 7.100 ;
        RECT 71.800 7.100 72.100 7.800 ;
        RECT 75.800 7.100 76.200 7.200 ;
        RECT 79.800 7.100 80.200 7.200 ;
        RECT 71.800 6.800 80.200 7.100 ;
        RECT 87.800 6.800 88.200 7.200 ;
        RECT 91.000 7.100 91.400 7.200 ;
        RECT 99.800 7.100 100.100 7.800 ;
        RECT 91.000 6.800 100.100 7.100 ;
        RECT 101.400 6.800 101.800 7.200 ;
        RECT 7.800 6.100 8.200 6.200 ;
        RECT 16.600 6.100 17.000 6.200 ;
        RECT 7.800 5.800 17.000 6.100 ;
        RECT 31.800 6.100 32.200 6.200 ;
        RECT 32.600 6.100 33.000 6.200 ;
        RECT 31.800 5.800 33.000 6.100 ;
        RECT 86.200 6.100 86.600 6.200 ;
        RECT 87.800 6.100 88.100 6.800 ;
        RECT 86.200 5.800 88.100 6.100 ;
        RECT 98.200 6.100 98.600 6.200 ;
        RECT 101.400 6.100 101.700 6.800 ;
        RECT 98.200 5.800 101.700 6.100 ;
        RECT 139.000 6.100 139.400 6.200 ;
        RECT 142.200 6.100 142.600 6.200 ;
        RECT 139.000 5.800 142.600 6.100 ;
        RECT 147.000 5.800 147.400 6.200 ;
        RECT 147.000 5.200 147.300 5.800 ;
        RECT 7.000 5.100 7.400 5.200 ;
        RECT 18.200 5.100 18.600 5.200 ;
        RECT 27.800 5.100 28.200 5.200 ;
        RECT 7.000 4.800 8.900 5.100 ;
        RECT 18.200 4.800 28.200 5.100 ;
        RECT 147.000 4.800 147.400 5.200 ;
        RECT 8.600 4.200 8.900 4.800 ;
        RECT 8.600 3.800 9.000 4.200 ;
      LAYER via3 ;
        RECT 87.000 126.800 87.400 127.200 ;
        RECT 135.000 126.800 135.400 127.200 ;
        RECT 35.000 124.800 35.400 125.200 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 127.000 124.800 127.400 125.200 ;
        RECT 40.600 121.800 41.000 122.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 147.000 121.800 147.400 122.200 ;
        RECT 145.400 116.800 145.800 117.200 ;
        RECT 41.400 114.800 41.800 115.200 ;
        RECT 126.200 114.800 126.600 115.200 ;
        RECT 86.200 113.800 86.600 114.200 ;
        RECT 41.400 109.800 41.800 110.200 ;
        RECT 43.800 109.800 44.200 110.200 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 147.000 105.800 147.400 106.200 ;
        RECT 90.200 104.800 90.600 105.200 ;
        RECT 107.000 104.800 107.400 105.200 ;
        RECT 146.200 104.800 146.600 105.200 ;
        RECT 104.600 99.800 105.000 100.200 ;
        RECT 147.000 96.800 147.400 97.200 ;
        RECT 11.000 95.800 11.400 96.200 ;
        RECT 61.400 94.800 61.800 95.200 ;
        RECT 107.000 93.800 107.400 94.200 ;
        RECT 68.600 91.800 69.000 92.200 ;
        RECT 147.800 89.800 148.200 90.200 ;
        RECT 145.400 88.800 145.800 89.200 ;
        RECT 95.800 86.800 96.200 87.200 ;
        RECT 107.000 86.800 107.400 87.200 ;
        RECT 132.600 86.800 133.000 87.200 ;
        RECT 105.400 83.800 105.800 84.200 ;
        RECT 149.400 83.800 149.800 84.200 ;
        RECT 91.800 82.800 92.200 83.200 ;
        RECT 94.200 80.800 94.600 81.200 ;
        RECT 139.800 79.800 140.200 80.200 ;
        RECT 59.000 76.800 59.400 77.200 ;
        RECT 64.600 76.800 65.000 77.200 ;
        RECT 139.800 76.800 140.200 77.200 ;
        RECT 143.800 75.800 144.200 76.200 ;
        RECT 139.000 74.800 139.400 75.200 ;
        RECT 87.800 71.800 88.200 72.200 ;
        RECT 30.200 70.800 30.600 71.200 ;
        RECT 40.600 70.800 41.000 71.200 ;
        RECT 146.200 68.800 146.600 69.200 ;
        RECT 11.000 66.800 11.400 67.200 ;
        RECT 124.600 66.800 125.000 67.200 ;
        RECT 99.800 65.800 100.200 66.200 ;
        RECT 15.800 64.800 16.200 65.200 ;
        RECT 76.600 64.800 77.000 65.200 ;
        RECT 119.800 64.800 120.200 65.200 ;
        RECT 130.200 64.800 130.600 65.200 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 103.000 53.800 103.400 54.200 ;
        RECT 80.600 52.800 81.000 53.200 ;
        RECT 20.600 51.800 21.000 52.200 ;
        RECT 85.400 51.800 85.800 52.200 ;
        RECT 95.800 51.800 96.200 52.200 ;
        RECT 104.600 51.800 105.000 52.200 ;
        RECT 91.800 50.800 92.200 51.200 ;
        RECT 93.400 50.800 93.800 51.200 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 147.000 48.800 147.400 49.200 ;
        RECT 38.200 47.800 38.600 48.200 ;
        RECT 98.200 47.800 98.600 48.200 ;
        RECT 117.400 46.800 117.800 47.200 ;
        RECT 96.600 45.800 97.000 46.200 ;
        RECT 87.800 42.800 88.200 43.200 ;
        RECT 86.200 41.800 86.600 42.200 ;
        RECT 137.400 41.800 137.800 42.200 ;
        RECT 65.400 40.800 65.800 41.200 ;
        RECT 27.800 38.800 28.200 39.200 ;
        RECT 82.200 32.800 82.600 33.200 ;
        RECT 90.200 30.800 90.600 31.200 ;
        RECT 151.000 29.800 151.400 30.200 ;
        RECT 89.400 28.800 89.800 29.200 ;
        RECT 15.800 22.800 16.200 23.200 ;
        RECT 126.200 15.800 126.600 16.200 ;
        RECT 84.600 14.800 85.000 15.200 ;
        RECT 47.800 12.800 48.200 13.200 ;
      LAYER metal4 ;
        RECT 87.000 126.800 87.400 127.200 ;
        RECT 135.000 126.800 135.400 127.200 ;
        RECT 147.800 126.800 148.200 127.200 ;
        RECT 87.000 126.200 87.300 126.800 ;
        RECT 87.000 125.800 87.400 126.200 ;
        RECT 112.600 126.100 113.000 126.200 ;
        RECT 113.400 126.100 113.800 126.200 ;
        RECT 112.600 125.800 113.800 126.100 ;
        RECT 135.000 125.200 135.300 126.800 ;
        RECT 35.000 124.800 35.400 125.200 ;
        RECT 127.000 125.100 127.400 125.200 ;
        RECT 126.200 124.800 127.400 125.100 ;
        RECT 135.000 124.800 135.400 125.200 ;
        RECT 35.000 107.200 35.300 124.800 ;
        RECT 40.600 121.800 41.000 122.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 35.000 106.800 35.400 107.200 ;
        RECT 11.000 95.800 11.400 96.200 ;
        RECT 11.000 67.200 11.300 95.800 ;
        RECT 29.400 94.100 29.800 94.200 ;
        RECT 29.400 93.800 30.500 94.100 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 17.400 68.800 17.800 69.200 ;
        RECT 11.000 66.800 11.400 67.200 ;
        RECT 15.800 64.800 16.200 65.200 ;
        RECT 15.800 23.200 16.100 64.800 ;
        RECT 17.400 42.200 17.700 68.800 ;
        RECT 20.600 52.200 20.900 73.800 ;
        RECT 30.200 71.200 30.500 93.800 ;
        RECT 40.600 71.200 40.900 121.800 ;
        RECT 41.400 114.800 41.800 115.200 ;
        RECT 41.400 112.200 41.700 114.800 ;
        RECT 41.400 111.800 41.800 112.200 ;
        RECT 41.400 110.200 41.700 111.800 ;
        RECT 41.400 109.800 41.800 110.200 ;
        RECT 43.800 109.800 44.200 110.200 ;
        RECT 43.800 95.200 44.100 109.800 ;
        RECT 61.400 105.800 61.800 106.200 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 61.400 95.200 61.700 105.800 ;
        RECT 64.600 101.800 65.000 102.200 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 61.400 94.800 61.800 95.200 ;
        RECT 47.800 90.800 48.200 91.200 ;
        RECT 30.200 70.800 30.600 71.200 ;
        RECT 40.600 70.800 41.000 71.200 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 20.600 51.800 21.000 52.200 ;
        RECT 17.400 41.800 17.800 42.200 ;
        RECT 27.800 39.200 28.100 54.800 ;
        RECT 38.200 48.100 38.600 48.200 ;
        RECT 39.000 48.100 39.400 48.200 ;
        RECT 38.200 47.800 39.400 48.100 ;
        RECT 43.800 48.100 44.200 48.200 ;
        RECT 44.600 48.100 45.000 48.200 ;
        RECT 43.800 47.800 45.000 48.100 ;
        RECT 27.800 38.800 28.200 39.200 ;
        RECT 15.800 22.800 16.200 23.200 ;
        RECT 47.800 13.200 48.100 90.800 ;
        RECT 58.200 81.800 58.600 82.200 ;
        RECT 58.200 69.200 58.500 81.800 ;
        RECT 59.000 76.800 59.400 77.200 ;
        RECT 59.000 75.200 59.300 76.800 ;
        RECT 59.000 74.800 59.400 75.200 ;
        RECT 58.200 68.800 58.600 69.200 ;
        RECT 51.000 59.800 51.400 60.200 ;
        RECT 51.000 29.200 51.300 59.800 ;
        RECT 59.000 54.200 59.300 74.800 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 59.000 49.200 59.300 53.800 ;
        RECT 59.000 48.800 59.400 49.200 ;
        RECT 61.400 46.200 61.700 94.800 ;
        RECT 64.600 84.200 64.900 101.800 ;
        RECT 68.600 92.200 68.900 105.800 ;
        RECT 68.600 91.800 69.000 92.200 ;
        RECT 74.200 84.200 74.500 121.800 ;
        RECT 126.200 115.200 126.500 124.800 ;
        RECT 147.000 121.800 147.400 122.200 ;
        RECT 145.400 116.800 145.800 117.200 ;
        RECT 126.200 114.800 126.600 115.200 ;
        RECT 86.200 114.100 86.600 114.200 ;
        RECT 85.400 113.800 86.600 114.100 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 85.400 90.200 85.700 113.800 ;
        RECT 119.800 113.200 120.100 113.800 ;
        RECT 87.800 112.800 88.200 113.200 ;
        RECT 119.800 112.800 120.200 113.200 ;
        RECT 85.400 89.800 85.800 90.200 ;
        RECT 82.200 86.800 82.600 87.200 ;
        RECT 64.600 83.800 65.000 84.200 ;
        RECT 74.200 83.800 74.600 84.200 ;
        RECT 64.600 77.100 65.000 77.200 ;
        RECT 63.800 76.800 65.000 77.100 ;
        RECT 63.800 67.200 64.100 76.800 ;
        RECT 76.600 67.800 77.000 68.200 ;
        RECT 63.800 66.800 64.200 67.200 ;
        RECT 76.600 65.200 76.900 67.800 ;
        RECT 76.600 64.800 77.000 65.200 ;
        RECT 65.400 56.800 65.800 57.200 ;
        RECT 61.400 45.800 61.800 46.200 ;
        RECT 65.400 41.200 65.700 56.800 ;
        RECT 80.600 52.800 81.000 53.200 ;
        RECT 65.400 40.800 65.800 41.200 ;
        RECT 80.600 38.200 80.900 52.800 ;
        RECT 80.600 37.800 81.000 38.200 ;
        RECT 82.200 33.200 82.500 86.800 ;
        RECT 87.800 72.200 88.100 112.800 ;
        RECT 119.800 109.200 120.100 112.800 ;
        RECT 139.800 109.800 140.200 110.200 ;
        RECT 119.800 108.800 120.200 109.200 ;
        RECT 97.400 107.800 97.800 108.200 ;
        RECT 90.200 104.800 90.600 105.200 ;
        RECT 88.600 95.800 89.000 96.200 ;
        RECT 88.600 80.200 88.900 95.800 ;
        RECT 90.200 85.200 90.500 104.800 ;
        RECT 94.200 93.800 94.600 94.200 ;
        RECT 90.200 84.800 90.600 85.200 ;
        RECT 88.600 79.800 89.000 80.200 ;
        RECT 89.400 78.800 89.800 79.200 ;
        RECT 87.800 71.800 88.200 72.200 ;
        RECT 88.600 67.100 89.000 67.200 ;
        RECT 89.400 67.100 89.700 78.800 ;
        RECT 88.600 66.800 89.700 67.100 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 85.400 51.800 85.800 52.200 ;
        RECT 85.400 36.200 85.700 51.800 ;
        RECT 88.600 48.200 88.900 54.800 ;
        RECT 86.200 47.800 86.600 48.200 ;
        RECT 88.600 47.800 89.000 48.200 ;
        RECT 86.200 42.200 86.500 47.800 ;
        RECT 87.800 42.800 88.200 43.200 ;
        RECT 86.200 41.800 86.600 42.200 ;
        RECT 87.800 37.200 88.100 42.800 ;
        RECT 87.800 36.800 88.200 37.200 ;
        RECT 85.400 35.800 85.800 36.200 ;
        RECT 82.200 32.800 82.600 33.200 ;
        RECT 84.600 29.800 85.000 30.200 ;
        RECT 51.000 28.800 51.400 29.200 ;
        RECT 84.600 15.200 84.900 29.800 ;
        RECT 87.800 25.200 88.100 36.800 ;
        RECT 89.400 29.200 89.700 66.800 ;
        RECT 90.200 74.200 90.500 84.800 ;
        RECT 91.800 82.800 92.200 83.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 90.200 31.200 90.500 73.800 ;
        RECT 91.800 68.200 92.100 82.800 ;
        RECT 94.200 81.200 94.500 93.800 ;
        RECT 95.800 87.100 96.200 87.200 ;
        RECT 96.600 87.100 97.000 87.200 ;
        RECT 95.800 86.800 97.000 87.100 ;
        RECT 97.400 86.100 97.700 107.800 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 98.200 94.200 98.500 106.800 ;
        RECT 107.000 104.800 107.400 105.200 ;
        RECT 104.600 102.800 105.000 103.200 ;
        RECT 104.600 100.200 104.900 102.800 ;
        RECT 104.600 99.800 105.000 100.200 ;
        RECT 105.400 99.800 105.800 100.200 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 96.600 85.800 97.700 86.100 ;
        RECT 94.200 80.800 94.600 81.200 ;
        RECT 93.400 73.800 93.800 74.200 ;
        RECT 91.800 67.800 92.200 68.200 ;
        RECT 91.800 52.800 92.200 53.200 ;
        RECT 91.800 51.200 92.100 52.800 ;
        RECT 93.400 51.200 93.700 73.800 ;
        RECT 95.800 53.800 96.200 54.200 ;
        RECT 95.800 52.200 96.100 53.800 ;
        RECT 95.800 51.800 96.200 52.200 ;
        RECT 91.800 50.800 92.200 51.200 ;
        RECT 93.400 50.800 93.800 51.200 ;
        RECT 96.600 46.200 96.900 85.800 ;
        RECT 105.400 84.200 105.700 99.800 ;
        RECT 107.000 94.200 107.300 104.800 ;
        RECT 123.800 103.100 124.200 103.200 ;
        RECT 124.600 103.100 125.000 103.200 ;
        RECT 123.800 102.800 125.000 103.100 ;
        RECT 107.000 93.800 107.400 94.200 ;
        RECT 107.000 87.200 107.300 93.800 ;
        RECT 107.000 86.800 107.400 87.200 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 132.600 87.100 133.000 87.200 ;
        RECT 131.800 86.800 133.000 87.100 ;
        RECT 139.000 85.800 139.400 86.200 ;
        RECT 105.400 83.800 105.800 84.200 ;
        RECT 124.600 77.800 125.000 78.200 ;
        RECT 135.000 77.800 135.400 78.200 ;
        RECT 124.600 67.200 124.900 77.800 ;
        RECT 124.600 66.800 125.000 67.200 ;
        RECT 99.800 65.800 100.200 66.200 ;
        RECT 99.800 65.200 100.100 65.800 ;
        RECT 124.600 65.200 124.900 66.800 ;
        RECT 99.800 64.800 100.200 65.200 ;
        RECT 119.000 65.100 119.400 65.200 ;
        RECT 119.800 65.100 120.200 65.200 ;
        RECT 119.000 64.800 120.200 65.100 ;
        RECT 124.600 64.800 125.000 65.200 ;
        RECT 129.400 65.100 129.800 65.200 ;
        RECT 130.200 65.100 130.600 65.200 ;
        RECT 129.400 64.800 130.600 65.100 ;
        RECT 135.000 56.200 135.300 77.800 ;
        RECT 139.000 75.200 139.300 85.800 ;
        RECT 139.800 80.200 140.100 109.800 ;
        RECT 145.400 95.200 145.700 116.800 ;
        RECT 146.200 112.800 146.600 113.200 ;
        RECT 146.200 105.200 146.500 112.800 ;
        RECT 147.000 106.200 147.300 121.800 ;
        RECT 147.000 105.800 147.400 106.200 ;
        RECT 146.200 104.800 146.600 105.200 ;
        RECT 147.000 96.800 147.400 97.200 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 145.400 88.800 145.800 89.200 ;
        RECT 144.600 86.800 145.000 87.200 ;
        RECT 139.800 79.800 140.200 80.200 ;
        RECT 139.800 77.200 140.100 79.800 ;
        RECT 139.800 76.800 140.200 77.200 ;
        RECT 139.800 75.200 140.100 76.800 ;
        RECT 143.800 75.800 144.200 76.200 ;
        RECT 139.000 74.800 139.400 75.200 ;
        RECT 139.800 74.800 140.200 75.200 ;
        RECT 137.400 73.800 137.800 74.200 ;
        RECT 137.400 67.200 137.700 73.800 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 135.000 55.800 135.400 56.200 ;
        RECT 98.200 54.100 98.600 54.200 ;
        RECT 97.400 53.800 98.600 54.100 ;
        RECT 102.200 54.100 102.600 54.200 ;
        RECT 103.000 54.100 103.400 54.200 ;
        RECT 102.200 53.800 103.400 54.100 ;
        RECT 97.400 49.200 97.700 53.800 ;
        RECT 103.000 50.200 103.300 53.800 ;
        RECT 137.400 53.200 137.700 66.800 ;
        RECT 137.400 53.100 137.800 53.200 ;
        RECT 138.200 53.100 138.600 53.200 ;
        RECT 137.400 52.800 138.600 53.100 ;
        RECT 104.600 51.800 105.000 52.200 ;
        RECT 131.000 51.800 131.400 52.200 ;
        RECT 103.000 49.800 103.400 50.200 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 98.200 47.800 98.600 48.200 ;
        RECT 98.200 46.200 98.500 47.800 ;
        RECT 104.600 47.200 104.900 51.800 ;
        RECT 104.600 46.800 105.000 47.200 ;
        RECT 116.600 47.100 117.000 47.200 ;
        RECT 117.400 47.100 117.800 47.200 ;
        RECT 116.600 46.800 117.800 47.100 ;
        RECT 96.600 45.800 97.000 46.200 ;
        RECT 98.200 45.800 98.600 46.200 ;
        RECT 125.400 31.800 125.800 32.200 ;
        RECT 90.200 30.800 90.600 31.200 ;
        RECT 89.400 28.800 89.800 29.200 ;
        RECT 87.800 24.800 88.200 25.200 ;
        RECT 125.400 16.100 125.700 31.800 ;
        RECT 131.000 27.200 131.300 51.800 ;
        RECT 137.400 47.800 137.800 48.200 ;
        RECT 137.400 42.200 137.700 47.800 ;
        RECT 137.400 41.800 137.800 42.200 ;
        RECT 131.000 26.800 131.400 27.200 ;
        RECT 143.800 26.200 144.100 75.800 ;
        RECT 144.600 45.200 144.900 86.800 ;
        RECT 145.400 84.200 145.700 88.800 ;
        RECT 145.400 83.800 145.800 84.200 ;
        RECT 145.400 76.800 145.800 77.200 ;
        RECT 144.600 44.800 145.000 45.200 ;
        RECT 143.800 25.800 144.200 26.200 ;
        RECT 145.400 25.200 145.700 76.800 ;
        RECT 147.000 74.200 147.300 96.800 ;
        RECT 147.800 94.200 148.100 126.800 ;
        RECT 148.600 114.800 149.000 115.200 ;
        RECT 147.800 93.800 148.200 94.200 ;
        RECT 147.800 89.800 148.200 90.200 ;
        RECT 147.000 73.800 147.400 74.200 ;
        RECT 146.200 68.800 146.600 69.200 ;
        RECT 146.200 54.200 146.500 68.800 ;
        RECT 147.800 56.200 148.100 89.800 ;
        RECT 147.800 55.800 148.200 56.200 ;
        RECT 146.200 53.800 146.600 54.200 ;
        RECT 147.000 48.800 147.400 49.200 ;
        RECT 146.200 35.800 146.600 36.200 ;
        RECT 145.400 24.800 145.800 25.200 ;
        RECT 146.200 19.200 146.500 35.800 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 126.200 16.100 126.600 16.200 ;
        RECT 125.400 15.800 126.600 16.100 ;
        RECT 84.600 14.800 85.000 15.200 ;
        RECT 47.800 12.800 48.200 13.200 ;
        RECT 147.000 5.200 147.300 48.800 ;
        RECT 148.600 17.200 148.900 114.800 ;
        RECT 149.400 108.800 149.800 109.200 ;
        RECT 149.400 84.200 149.700 108.800 ;
        RECT 150.200 95.800 150.600 96.200 ;
        RECT 149.400 83.800 149.800 84.200 ;
        RECT 150.200 73.200 150.500 95.800 ;
        RECT 151.000 88.800 151.400 89.200 ;
        RECT 150.200 72.800 150.600 73.200 ;
        RECT 151.000 30.200 151.300 88.800 ;
        RECT 151.000 29.800 151.400 30.200 ;
        RECT 148.600 16.800 149.000 17.200 ;
        RECT 147.000 4.800 147.400 5.200 ;
      LAYER via4 ;
        RECT 39.000 47.800 39.400 48.200 ;
        RECT 96.600 86.800 97.000 87.200 ;
        RECT 124.600 102.800 125.000 103.200 ;
        RECT 138.200 52.800 138.600 53.200 ;
      LAYER metal5 ;
        RECT 87.000 126.100 87.400 126.200 ;
        RECT 112.600 126.100 113.000 126.200 ;
        RECT 87.000 125.800 113.000 126.100 ;
        RECT 87.800 113.100 88.200 113.200 ;
        RECT 119.800 113.100 120.200 113.200 ;
        RECT 87.800 112.800 120.200 113.100 ;
        RECT 104.600 103.100 105.000 103.200 ;
        RECT 124.600 103.100 125.000 103.200 ;
        RECT 104.600 102.800 125.000 103.100 ;
        RECT 96.600 87.100 97.000 87.200 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 96.600 86.800 132.200 87.100 ;
        RECT 99.800 65.100 100.200 65.200 ;
        RECT 119.000 65.100 119.400 65.200 ;
        RECT 129.400 65.100 129.800 65.200 ;
        RECT 99.800 64.800 129.800 65.100 ;
        RECT 95.800 54.100 96.200 54.200 ;
        RECT 102.200 54.100 102.600 54.200 ;
        RECT 95.800 53.800 102.600 54.100 ;
        RECT 91.800 53.100 92.200 53.200 ;
        RECT 138.200 53.100 138.600 53.200 ;
        RECT 91.800 52.800 138.600 53.100 ;
        RECT 39.000 48.100 39.400 48.200 ;
        RECT 43.800 48.100 44.200 48.200 ;
        RECT 39.000 47.800 44.200 48.100 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 116.600 47.100 117.000 47.200 ;
        RECT 104.600 46.800 117.000 47.100 ;
  END
END pipeline
END LIBRARY

