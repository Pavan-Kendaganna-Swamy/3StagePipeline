* NGSPICE file created from pipeline.ext - technology: scmos

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt pipeline vdd gnd A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3]
+ B[4] B[5] B[6] B[7] C[0] C[1] C[2] C[3] C[4] C[5] C[6] C[7] D[0] D[1] D[2] D[3]
+ D[4] D[5] D[6] D[7] clk F[0] F[1] F[2] F[3] F[4] F[5] F[6] F[7]
XAND2X2_5 OR2X2_3/Y AND2X2_5/B gnd INVX1_37/A vdd AND2X2
XNAND2X1_32 OAI21X1_31/Y OAI21X1_30/Y gnd OAI21X1_40/B vdd NAND2X1
XNAND2X1_43 NAND2X1_43/A NAND2X1_43/B gnd NAND2X1_43/Y vdd NAND2X1
XNAND2X1_54 AND2X2_6/Y XOR2X1_19/A gnd NAND2X1_54/Y vdd NAND2X1
XNAND2X1_10 AOI22X1_3/A INVX2_1/A gnd NOR2X1_9/B vdd NAND2X1
XNAND2X1_21 BUFX4_8/Y INVX1_15/A gnd OAI22X1_5/A vdd NAND2X1
XOAI22X1_3 NOR2X1_7/B NOR2X1_13/A AOI22X1_4/Y INVX2_4/A gnd OAI22X1_3/Y vdd OAI22X1
XFILL_11_1_0 gnd vdd FILL
XOAI21X1_19 AOI21X1_11/Y OAI21X1_16/B INVX1_10/Y gnd NAND2X1_23/B vdd OAI21X1
XXNOR2X1_6 NOR3X1_5/A INVX2_6/Y gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_8_1_0 gnd vdd FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_44 AND2X2_2/Y XOR2X1_6/A gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_55 XOR2X1_21/A XOR2X1_21/B gnd NAND2X1_55/Y vdd NAND2X1
XNAND2X1_33 NAND2X1_33/A INVX4_1/A gnd XNOR2X1_4/B vdd NAND2X1
XAOI22X1_1 BUFX4_8/Y AOI22X1_3/B BUFX4_4/Y NAND2X1_3/B gnd INVX1_9/A vdd AOI22X1
XNAND2X1_11 BUFX4_1/Y AOI22X1_3/B gnd NOR2X1_7/A vdd NAND2X1
XNAND2X1_22 NOR2X1_7/A NOR2X1_7/B gnd AOI21X1_15/B vdd NAND2X1
XOAI22X1_4 OAI22X1_4/A XOR2X1_3/A AOI22X1_3/Y INVX1_12/A gnd XOR2X1_4/B vdd OAI22X1
XFILL_11_1_1 gnd vdd FILL
XXNOR2X1_7 NOR3X1_5/A INVX2_6/A gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XNAND2X1_56 INVX1_44/A XNOR2X1_25/A gnd OAI21X1_58/C vdd NAND2X1
XNAND2X1_45 B[4] A[4] gnd NAND2X1_47/A vdd NAND2X1
XNAND2X1_23 NAND3X1_18/Y NAND2X1_23/B gnd OAI21X1_23/B vdd NAND2X1
XNAND2X1_12 INVX1_2/A NAND2X1_3/B gnd INVX2_3/A vdd NAND2X1
XAOI22X1_2 BUFX4_7/Y AOI22X1_4/D INVX1_4/A AOI22X1_3/B gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_34 NAND2X1_34/A NAND2X1_3/B gnd INVX2_6/A vdd NAND2X1
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B OAI22X1_5/C INVX1_13/A gnd NOR3X1_4/A vdd OAI22X1
XXNOR2X1_8 NOR3X1_4/A INVX2_6/Y gnd XNOR2X1_8/Y vdd XNOR2X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_9_1 gnd vdd FILL
XAND2X2_8 INVX1_49/Y AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XAOI22X1_3 AOI22X1_3/A AOI22X1_3/B INVX1_7/A NAND2X1_3/B gnd AOI22X1_3/Y vdd AOI22X1
XNAND2X1_46 XOR2X1_9/B XOR2X1_9/A gnd NAND2X1_47/B vdd NAND2X1
XNAND2X1_57 NOR2X1_38/A NOR2X1_38/B gnd INVX1_45/A vdd NAND2X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR2X1_8/Y gnd NOR3X1_1/Y vdd NOR3X1
XNAND2X1_24 INVX1_7/A NAND2X1_3/B gnd AOI21X1_24/C vdd NAND2X1
XNAND2X1_13 BUFX4_5/Y AOI22X1_4/D gnd NOR2X1_7/B vdd NAND2X1
XNAND2X1_35 AOI22X1_3/A AOI22X1_4/D gnd XOR2X1_3/B vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XXNOR2X1_9 NOR3X1_4/A INVX2_6/A gnd XNOR2X1_9/Y vdd XNOR2X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_9_2 gnd vdd FILL
XAND2X2_9 INVX1_1/Y AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XXOR2X1_20 XOR2X1_20/A XOR2X1_20/B gnd XOR2X1_20/Y vdd XOR2X1
XAOI22X1_4 BUFX4_7/Y INVX1_15/A BUFX4_4/Y AOI22X1_4/D gnd AOI22X1_4/Y vdd AOI22X1
XNAND2X1_58 NOR2X1_40/A NOR2X1_40/B gnd INVX1_46/A vdd NAND2X1
XNAND2X1_47 NAND2X1_47/A NAND2X1_47/B gnd XOR2X1_10/A vdd NAND2X1
XNAND2X1_36 BUFX4_4/Y AOI22X1_5/B gnd OAI22X1_5/B vdd NAND2X1
XNOR3X1_2 NOR3X1_2/A OR2X2_1/Y NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XNAND2X1_14 NAND3X1_7/Y OAI21X1_13/Y gnd OR2X2_1/A vdd NAND2X1
XNAND2X1_25 NAND2X1_34/A INVX2_1/A gnd INVX1_12/A vdd NAND2X1
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XFILL_3_0_1 gnd vdd FILL
XXOR2X1_21 XOR2X1_21/A XOR2X1_21/B gnd INVX1_41/A vdd XOR2X1
XXOR2X1_10 XOR2X1_10/A NOR2X1_27/Y gnd XOR2X1_10/Y vdd XOR2X1
XNAND2X1_37 INVX1_2/A INVX1_15/A gnd INVX1_17/A vdd NAND2X1
XAOI22X1_5 BUFX4_8/Y AOI22X1_5/B INVX1_4/A INVX1_15/A gnd OAI22X1_5/C vdd AOI22X1
XNAND2X1_48 B[6] A[6] gnd NAND2X1_48/Y vdd NAND2X1
XNAND2X1_59 NOR2X1_42/A NOR2X1_42/B gnd INVX1_47/A vdd NAND2X1
XNAND2X1_15 INVX1_7/A INVX4_1/A gnd NOR2X1_9/A vdd NAND2X1
XNAND2X1_26 AOI22X1_3/A AOI22X1_3/B gnd NAND2X1_26/Y vdd NAND2X1
XNOR3X1_3 NOR3X1_3/A INVX1_17/A NOR3X1_3/C gnd NOR3X1_4/C vdd NOR3X1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XXOR2X1_11 XOR2X1_11/A XOR2X1_11/B gnd XOR2X1_11/Y vdd XOR2X1
XXOR2X1_22 XOR2X1_22/A XOR2X1_22/B gnd XOR2X1_22/Y vdd XOR2X1
XFILL_1_1_0 gnd vdd FILL
XNAND3X1_1 OAI21X1_3/Y INVX1_6/Y NAND3X1_1/C gnd NAND3X1_3/B vdd NAND3X1
XNAND2X1_38 NAND3X1_54/A BUFX4_6/Y gnd NAND2X1_38/Y vdd NAND2X1
XNAND2X1_49 XOR2X1_13/B XOR2X1_13/A gnd NAND2X1_49/Y vdd NAND2X1
XAOI22X1_6 NOR2X1_14/Y NOR2X1_8/Y OR2X2_2/A AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XNAND2X1_16 NAND2X1_34/A INVX4_1/A gnd INVX1_10/A vdd NAND2X1
XNAND2X1_27 INVX1_7/A AOI22X1_3/B gnd XOR2X1_3/A vdd NAND2X1
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XXOR2X1_12 C[0] D[0] gnd XOR2X1_12/Y vdd XOR2X1
XNAND3X1_2 INVX1_6/A OAI21X1_5/Y OAI21X1_4/Y gnd NAND3X1_3/C vdd NAND3X1
XNAND2X1_28 OAI21X1_25/Y OAI21X1_24/Y gnd AOI21X1_39/A vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XNAND2X1_39 XOR2X1_1/B XOR2X1_1/A gnd INVX2_7/A vdd NAND2X1
XNAND2X1_17 AOI22X1_3/A NAND2X1_3/B gnd OAI22X1_4/A vdd NAND2X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_5/Y vdd NOR3X1
XXOR2X1_2 XOR2X1_4/B XOR2X1_2/B gnd XOR2X1_2/Y vdd XOR2X1
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_13 XOR2X1_13/A XOR2X1_13/B gnd XOR2X1_13/Y vdd XOR2X1
XNAND3X1_3 INVX1_5/Y NAND3X1_3/B NAND3X1_3/C gnd NAND3X1_3/Y vdd NAND3X1
XNAND2X1_29 INVX1_4/A INVX1_15/A gnd NOR2X1_13/A vdd NAND2X1
XNAND2X1_18 NAND3X1_10/Y OAI21X1_16/Y gnd AOI21X1_29/A vdd NAND2X1
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd XOR2X1_3/Y vdd XOR2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_12_0_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XBUFX4_1 BUFX4_4/A gnd BUFX4_1/Y vdd BUFX4
XFILL_4_1_0 gnd vdd FILL
XXOR2X1_14 XOR2X1_14/A XOR2X1_14/B gnd XOR2X1_14/Y vdd XOR2X1
XNAND3X1_4 NOR2X1_3/Y NAND3X1_3/Y OAI21X1_6/Y gnd NOR3X1_1/A vdd NAND3X1
XNAND2X1_19 BUFX4_4/Y AOI22X1_4/D gnd NOR2X1_12/A vdd NAND2X1
XFILL_5_1 gnd vdd FILL
XAOI21X1_50 XOR2X1_7/B XOR2X1_7/A AND2X2_3/Y gnd AOI21X1_50/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XOAI21X1_1 INVX1_4/Y INVX2_1/Y OAI22X1_1/A gnd OAI21X1_1/Y vdd OAI21X1
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XXOR2X1_15 C[6] D[6] gnd XOR2X1_16/B vdd XOR2X1
XFILL_4_1_1 gnd vdd FILL
XBUFX4_2 BUFX4_4/A gnd BUFX4_2/Y vdd BUFX4
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 NAND3X1_5/A AOI21X1_9/A OAI21X1_9/Y gnd NAND3X1_7/B vdd NAND3X1
XAOI21X1_40 AOI21X1_45/A AOI21X1_45/B XOR2X1_4/A gnd OAI21X1_41/A vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_2 NOR2X1_4/A NOR2X1_5/A OAI21X1_1/Y gnd XNOR2X1_1/A vdd OAI21X1
XAOI21X1_51 INVX1_29/Y XOR2X1_10/A NOR2X1_25/Y gnd XOR2X1_11/A vdd AOI21X1
XXOR2X1_5 B[1] A[1] gnd XOR2X1_6/A vdd XOR2X1
XDFFPOSX1_40 NAND2X1_3/B CLKBUF1_6/Y XOR2X1_20/Y gnd vdd DFFPOSX1
XXOR2X1_16 XOR2X1_16/A XOR2X1_16/B gnd XOR2X1_16/Y vdd XOR2X1
XBUFX4_3 BUFX4_4/A gnd INVX1_4/A vdd BUFX4
XNAND3X1_6 NAND3X1_6/A AOI21X1_8/C NAND3X1_6/C gnd NAND3X1_6/Y vdd NAND3X1
XAOI21X1_41 AOI21X1_36/A AOI21X1_36/B XOR2X1_3/Y gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_30 NAND3X1_46/A NAND3X1_42/Y NAND3X1_45/B gnd AOI21X1_33/C vdd AOI21X1
XAOI21X1_52 INVX2_8/A XNOR2X1_21/A INVX1_35/A gnd AOI21X1_52/Y vdd AOI21X1
XOAI21X1_3 NOR2X1_5/Y INVX1_9/A INVX2_2/A gnd OAI21X1_3/Y vdd OAI21X1
XFILL_10_1_0 gnd vdd FILL
XXOR2X1_6 XOR2X1_6/A AND2X2_2/Y gnd XOR2X1_6/Y vdd XOR2X1
XDFFPOSX1_41 AOI22X1_3/B CLKBUF1_4/Y XNOR2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 AND2X2_6/B CLKBUF1_5/Y XOR2X1_12/Y gnd vdd DFFPOSX1
XFILL_7_1_0 gnd vdd FILL
XBUFX4_4 BUFX4_4/A gnd BUFX4_4/Y vdd BUFX4
XXOR2X1_17 C[7] D[7] gnd XOR2X1_17/Y vdd XOR2X1
XNAND3X1_7 INVX1_8/Y NAND3X1_7/B NAND3X1_6/Y gnd NAND3X1_7/Y vdd NAND3X1
XBUFX2_1 BUFX2_1/A gnd F[0] vdd BUFX2
XAOI21X1_1 INVX1_3/A OAI21X1_1/Y NOR2X1_4/Y gnd INVX1_6/A vdd AOI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XXNOR2X1_20 C[3] D[3] gnd XOR2X1_14/B vdd XNOR2X1
XAOI21X1_42 NAND3X1_37/B NAND3X1_37/C OAI22X1_3/Y gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_31 NAND3X1_36/Y AOI21X1_31/B AOI21X1_31/C gnd AOI21X1_31/Y vdd AOI21X1
XOAI21X1_4 INVX1_2/Y INVX2_1/Y NOR2X1_6/Y gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_20 NAND3X1_25/Y OAI21X1_32/C INVX2_5/A gnd NOR3X1_2/C vdd AOI21X1
XAOI21X1_53 NOR2X1_32/Y XNOR2X1_21/A AOI21X1_53/C gnd XOR2X1_16/A vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B gnd XOR2X1_7/Y vdd XOR2X1
XFILL_10_1_1 gnd vdd FILL
XDFFPOSX1_42 AOI22X1_4/D CLKBUF1_4/Y XNOR2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX1_40/A CLKBUF1_5/Y XNOR2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 INVX1_11/A CLKBUF1_1/Y DFFPOSX1_12/Q gnd vdd DFFPOSX1
XFILL_7_1_1 gnd vdd FILL
XXOR2X1_18 INVX1_39/A INVX1_40/A gnd XOR2X1_19/A vdd XOR2X1
XBUFX4_5 BUFX4_7/A gnd BUFX4_5/Y vdd BUFX4
XBUFX2_2 BUFX2_2/A gnd F[1] vdd BUFX2
XNAND3X1_8 AOI22X1_3/A NAND2X1_3/B NAND3X1_8/C gnd NAND3X1_8/Y vdd NAND3X1
XXNOR2X1_10 XOR2X1_2/B XNOR2X1_4/B gnd INVX1_19/A vdd XNOR2X1
XAOI21X1_2 OAI21X1_5/Y OAI21X1_4/Y INVX1_6/A gnd AOI21X1_4/C vdd AOI21X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XXNOR2X1_21 XNOR2X1_21/A INVX2_8/Y gnd XNOR2X1_21/Y vdd XNOR2X1
XAOI21X1_43 AOI21X1_46/A AOI21X1_46/B AOI21X1_43/C gnd OAI21X1_41/B vdd AOI21X1
XAOI21X1_10 NAND3X1_7/Y OAI21X1_13/Y OAI21X1_14/Y gnd NOR3X1_1/B vdd AOI21X1
XAOI21X1_32 NAND3X1_48/Y NAND3X1_50/Y NAND3X1_72/B gnd NOR2X1_15/A vdd AOI21X1
XAOI21X1_54 XOR2X1_20/B XOR2X1_20/A AND2X2_7/Y gnd XNOR2X1_24/A vdd AOI21X1
XOAI21X1_5 NOR2X1_5/Y INVX1_9/A INVX2_2/Y gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_21 INVX2_5/A NAND3X1_25/Y AOI21X1_17/Y gnd NAND3X1_48/C vdd AOI21X1
XFILL_3_2 gnd vdd FILL
XXOR2X1_8 B[4] A[4] gnd XOR2X1_9/B vdd XOR2X1
XDFFPOSX1_43 INVX1_15/A CLKBUF1_4/Y NOR2X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 NAND2X1_33/A CLKBUF1_1/Y DFFPOSX1_13/Q gnd vdd DFFPOSX1
XDFFPOSX1_32 AND2X2_7/B CLKBUF1_5/Y XOR2X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 DFFPOSX1_10/Q CLKBUF1_6/Y D[4] gnd vdd DFFPOSX1
XXOR2X1_19 XOR2X1_19/A AND2X2_6/Y gnd XOR2X1_19/Y vdd XOR2X1
XBUFX4_6 BUFX4_7/A gnd BUFX4_6/Y vdd BUFX4
XBUFX2_3 BUFX2_3/A gnd F[2] vdd BUFX2
XNAND3X1_9 INVX1_7/A INVX2_1/A OAI22X1_4/A gnd NAND3X1_9/Y vdd NAND3X1
XAOI21X1_3 OAI21X1_3/Y NAND3X1_1/C INVX1_6/Y gnd OAI21X1_6/B vdd AOI21X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XXNOR2X1_11 XOR2X1_4/A XOR2X1_4/B gnd NAND3X1_66/C vdd XNOR2X1
XXNOR2X1_22 AOI21X1_52/Y INVX1_37/A gnd XNOR2X1_22/Y vdd XNOR2X1
XNOR2X1_1 NOR2X1_4/A NOR2X1_1/B gnd INVX1_1/A vdd NOR2X1
XAOI21X1_33 XOR2X1_1/Y AOI21X1_33/B AOI21X1_33/C gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_55 INVX1_45/A INVX1_46/A INVX1_48/Y gnd INVX1_49/A vdd AOI21X1
XOAI21X1_6 AOI21X1_4/C OAI21X1_6/B INVX1_5/A gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_11 INVX1_7/A INVX2_1/A OAI22X1_4/A gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_22 NAND3X1_14/B OAI21X1_17/Y OAI22X1_2/Y gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_44 NAND3X1_63/Y OAI21X1_41/Y AOI21X1_33/Y gnd NOR2X1_17/A vdd AOI21X1
XXOR2X1_9 XOR2X1_9/A XOR2X1_9/B gnd XOR2X1_9/Y vdd XOR2X1
XDFFPOSX1_11 DFFPOSX1_11/Q CLKBUF1_6/Y D[5] gnd vdd DFFPOSX1
XDFFPOSX1_44 AOI22X1_5/B CLKBUF1_4/Y AND2X2_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 XOR2X1_21/B CLKBUF1_2/Y XOR2X1_14/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_22 BUFX2_1/A CLKBUF1_3/Y NOR2X1_19/Y gnd vdd DFFPOSX1
XFILL_13_1 gnd vdd FILL
XBUFX4_7 BUFX4_7/A gnd BUFX4_7/Y vdd BUFX4
XBUFX2_4 BUFX2_4/A gnd F[3] vdd BUFX2
XAOI21X1_4 INVX1_5/Y NAND3X1_3/C AOI21X1_4/C gnd OR2X2_1/B vdd AOI21X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XNOR2X1_2 INVX1_2/Y INVX4_1/Y gnd INVX1_3/A vdd NOR2X1
XXNOR2X1_23 XNOR2X1_23/A XOR2X1_17/Y gnd XNOR2X1_23/Y vdd XNOR2X1
XXNOR2X1_12 OR2X2_2/A INVX2_7/A gnd NAND2X1_40/B vdd XNOR2X1
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B INVX1_19/Y gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_34 BUFX4_2/Y AOI22X1_5/B NAND2X1_38/Y gnd NOR3X1_3/A vdd AOI21X1
XAOI21X1_56 NAND3X1_3/Y OAI21X1_6/Y NOR2X1_3/Y gnd NOR2X1_47/A vdd AOI21X1
XOAI21X1_7 INVX1_7/Y INVX4_1/Y NOR2X1_9/B gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_12 AOI22X1_3/A NAND2X1_3/B NAND3X1_8/C gnd OAI21X1_16/B vdd AOI21X1
XAOI21X1_23 INVX1_7/A NAND2X1_3/B NAND2X1_26/Y gnd OAI21X1_30/A vdd AOI21X1
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_34 INVX1_43/A CLKBUF1_2/Y XNOR2X1_21/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_23 BUFX2_2/A CLKBUF1_3/Y AND2X2_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 DFFPOSX1_12/Q CLKBUF1_5/Y D[6] gnd vdd DFFPOSX1
XDFFPOSX1_45 NAND3X1_54/A CLKBUF1_6/Y XOR2X1_22/Y gnd vdd DFFPOSX1
XFILL_13_2 gnd vdd FILL
XBUFX4_8 BUFX4_7/A gnd BUFX4_8/Y vdd BUFX4
XBUFX2_5 BUFX2_5/A gnd F[4] vdd BUFX2
XXNOR2X1_13 AOI21X1_50/Y NOR2X1_24/Y gnd DFFPOSX1_1/D vdd XNOR2X1
XXNOR2X1_24 XNOR2X1_24/A INVX1_41/A gnd XNOR2X1_24/Y vdd XNOR2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XAOI21X1_5 BUFX4_2/Y AOI22X1_3/B NOR2X1_7/B gnd AOI21X1_5/Y vdd AOI21X1
XAOI21X1_46 AOI21X1_46/A AOI21X1_46/B INVX1_19/A gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_57 NAND3X1_72/B OAI21X1_21/Y NOR3X1_1/Y gnd NOR2X1_48/A vdd AOI21X1
XNOR2X1_3 INVX1_1/Y NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_24 AOI22X1_3/A AOI22X1_3/B AOI21X1_24/C gnd OAI21X1_30/B vdd AOI21X1
XAOI21X1_35 NAND3X1_54/A BUFX4_7/Y OAI22X1_5/B gnd NOR3X1_3/C vdd AOI21X1
XAOI21X1_13 BUFX4_1/Y AOI22X1_4/D OAI22X1_5/A gnd OAI21X1_17/A vdd AOI21X1
XOAI21X1_8 INVX1_5/A NAND3X1_8/C OAI21X1_7/Y gnd INVX1_8/A vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XDFFPOSX1_46 AND2X2_6/A CLKBUF1_4/Y NOR2X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 NOR2X1_38/B CLKBUF1_2/Y XNOR2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 BUFX2_3/A CLKBUF1_3/Y AND2X2_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 DFFPOSX1_13/Q CLKBUF1_5/Y D[7] gnd vdd DFFPOSX1
XFILL_13_3 gnd vdd FILL
XBUFX2_6 BUFX2_6/A gnd F[5] vdd BUFX2
XNAND2X1_1 BUFX4_5/Y INVX2_1/A gnd NOR2X1_4/A vdd NAND2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XXNOR2X1_25 XNOR2X1_25/A INVX1_44/Y gnd XNOR2X1_25/Y vdd XNOR2X1
XDFFPOSX1_1 XOR2X1_21/A CLKBUF1_2/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XFILL_0_1_0 gnd vdd FILL
XXNOR2X1_14 B[6] A[6] gnd XOR2X1_11/B vdd XNOR2X1
XAOI21X1_6 BUFX4_6/Y AOI22X1_4/D NOR2X1_7/A gnd AOI21X1_6/Y vdd AOI21X1
XNOR2X1_4 NOR2X1_4/A NOR2X1_5/A gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_36 AOI21X1_36/A AOI21X1_36/B INVX1_16/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_47 OAI21X1_43/Y NAND3X1_66/Y AOI21X1_47/C gnd NOR2X1_17/B vdd AOI21X1
XAOI21X1_25 BUFX4_1/Y INVX1_15/A NOR2X1_13/B gnd OAI21X1_26/A vdd AOI21X1
XOAI21X1_9 AOI21X1_5/Y AOI21X1_6/Y INVX2_3/Y gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_14 BUFX4_5/Y INVX1_15/A NOR2X1_12/A gnd OAI21X1_17/B vdd AOI21X1
XFILL_1_3 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_25 BUFX2_4/A CLKBUF1_3/Y NOR2X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 NOR2X1_42/B CLKBUF1_5/Y XOR2X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 BUFX4_7/A CLKBUF1_1/Y DFFPOSX1_6/Q gnd vdd DFFPOSX1
XDFFPOSX1_47 INVX1_39/A CLKBUF1_6/Y XOR2X1_6/Y gnd vdd DFFPOSX1
XBUFX2_7 BUFX2_7/A gnd F[6] vdd BUFX2
XFILL_0_1_1 gnd vdd FILL
XINVX1_50 NOR2X1_3/Y gnd INVX1_50/Y vdd INVX1
XNAND2X1_2 BUFX4_1/Y INVX4_1/A gnd NOR2X1_1/B vdd NAND2X1
XAOI21X1_7 INVX2_2/Y INVX1_9/Y NOR2X1_5/Y gnd AOI21X1_8/C vdd AOI21X1
XXNOR2X1_26 DFFPOSX1_5/Q XNOR2X1_26/B gnd XOR2X1_22/B vdd XNOR2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XXNOR2X1_15 B[7] A[7] gnd XNOR2X1_16/B vdd XNOR2X1
XDFFPOSX1_2 INVX1_42/A CLKBUF1_4/Y XOR2X1_9/Y gnd vdd DFFPOSX1
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_37 AOI21X1_37/A AOI21X1_37/B INVX1_17/Y gnd NOR3X1_4/B vdd AOI21X1
XAOI21X1_26 BUFX4_5/Y AOI22X1_5/B NOR2X1_13/A gnd OAI21X1_26/B vdd AOI21X1
XAOI21X1_48 AOI21X1_48/A OAI21X1_45/Y AND2X2_11/A gnd NOR2X1_48/B vdd AOI21X1
XAOI21X1_15 INVX2_3/Y AOI21X1_15/B NOR2X1_7/Y gnd NAND3X1_19/A vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_48 AND2X2_7/A CLKBUF1_4/Y XOR2X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_37 XNOR2X1_26/B CLKBUF1_5/Y XNOR2X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 BUFX2_5/A CLKBUF1_3/Y AND2X2_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 BUFX4_4/A CLKBUF1_1/Y DFFPOSX1_7/Q gnd vdd DFFPOSX1
XBUFX2_8 BUFX2_8/A gnd F[7] vdd BUFX2
XNAND3X1_70 OR2X2_1/Y INVX1_21/Y INVX1_20/Y gnd AND2X2_11/A vdd NAND3X1
XNAND2X1_3 BUFX4_2/Y NAND2X1_3/B gnd NOR2X1_5/A vdd NAND2X1
XAOI21X1_8 NAND3X1_6/A NAND3X1_6/C AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XNOR2X1_6 INVX1_9/A NOR2X1_5/Y gnd NOR2X1_6/Y vdd NOR2X1
XXNOR2X1_16 XNOR2X1_16/A XNOR2X1_16/B gnd XNOR2X1_16/Y vdd XNOR2X1
XDFFPOSX1_3 NOR2X1_38/A CLKBUF1_2/Y XOR2X1_10/Y gnd vdd DFFPOSX1
XAOI21X1_38 AOI21X1_38/A AOI21X1_38/B AOI21X1_38/C gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_27 INVX2_4/Y OAI21X1_27/Y NOR2X1_12/Y gnd AOI21X1_38/C vdd AOI21X1
XAOI21X1_49 NAND3X1_72/Y NOR2X1_48/B NOR2X1_15/A gnd AOI21X1_49/Y vdd AOI21X1
XAOI21X1_16 INVX1_8/Y NAND3X1_6/Y AOI21X1_8/Y gnd NAND3X1_28/C vdd AOI21X1
XDFFPOSX1_16 INVX1_2/A CLKBUF1_1/Y DFFPOSX1_8/Q gnd vdd DFFPOSX1
XDFFPOSX1_27 BUFX2_6/A CLKBUF1_3/Y NOR2X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 INVX4_1/A CLKBUF1_1/Y NOR2X1_46/Y gnd vdd DFFPOSX1
XFILL_3_1_0 gnd vdd FILL
XNAND3X1_60 XNOR2X1_8/Y NAND3X1_59/Y NAND3X1_60/C gnd AOI21X1_46/A vdd NAND3X1
XFILL_11_0_0 gnd vdd FILL
XNAND3X1_71 NAND3X1_27/B OR2X2_1/Y OAI21X1_20/Y gnd AOI21X1_48/A vdd NAND3X1
XNAND2X1_4 BUFX4_6/Y NAND2X1_3/B gnd OAI22X1_1/A vdd NAND2X1
XAOI21X1_9 AOI21X1_9/A OAI21X1_9/Y NAND3X1_5/A gnd AOI21X1_9/Y vdd AOI21X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XINVX1_30 D[0] gnd INVX1_30/Y vdd INVX1
XXNOR2X1_17 C[1] D[1] gnd XNOR2X1_18/A vdd XNOR2X1
XDFFPOSX1_4 NOR2X1_42/A CLKBUF1_2/Y XOR2X1_11/Y gnd vdd DFFPOSX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XAOI21X1_39 AOI21X1_39/A AOI21X1_39/B AOI21X1_38/Y gnd XOR2X1_4/A vdd AOI21X1
XAOI21X1_17 NAND3X1_23/Y NAND3X1_24/Y NAND3X1_28/C gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 NAND3X1_15/Y OAI21X1_18/Y NAND3X1_19/A gnd AOI21X1_28/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XDFFPOSX1_28 BUFX2_7/A CLKBUF1_3/Y XNOR2X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_39 INVX2_1/A CLKBUF1_4/Y XOR2X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_17 AOI22X1_3/A CLKBUF1_6/Y DFFPOSX1_9/Q gnd vdd DFFPOSX1
XFILL_3_1_1 gnd vdd FILL
XNAND3X1_61 AOI21X1_46/A AOI21X1_43/C AOI21X1_46/B gnd NAND3X1_61/Y vdd NAND3X1
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_72 NAND3X1_48/Y NAND3X1_72/B NAND3X1_50/Y gnd NAND3X1_72/Y vdd NAND3X1
XNAND3X1_50 NAND3X1_49/Y NAND3X1_51/B OAI21X1_33/Y gnd NAND3X1_50/Y vdd NAND3X1
XNAND2X1_5 AOI22X1_3/A INVX4_1/A gnd INVX1_5/A vdd NAND2X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_20 NOR3X1_1/A gnd INVX1_20/Y vdd INVX1
XXNOR2X1_18 XNOR2X1_18/A NOR2X1_30/Y gnd XNOR2X1_18/Y vdd XNOR2X1
XINVX1_31 C[1] gnd INVX1_31/Y vdd INVX1
XDFFPOSX1_5 DFFPOSX1_5/Q CLKBUF1_2/Y XNOR2X1_16/Y gnd vdd DFFPOSX1
XNOR2X1_8 OR2X2_1/B OR2X2_1/A gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 NAND3X1_17/Y NAND3X1_21/Y AOI21X1_18/C gnd OAI21X1_32/A vdd AOI21X1
XAOI21X1_29 AOI21X1_29/A NAND3X1_16/Y AOI21X1_28/Y gnd NAND3X1_45/B vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XDFFPOSX1_29 BUFX2_8/A CLKBUF1_3/Y NAND2X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_18 INVX1_7/A CLKBUF1_6/Y DFFPOSX1_10/Q gnd vdd DFFPOSX1
XNAND3X1_62 XOR2X1_4/A AOI21X1_45/A AOI21X1_45/B gnd NAND3X1_62/Y vdd NAND3X1
XNAND3X1_40 NAND3X1_36/Y AOI21X1_31/B AOI21X1_31/C gnd NAND3X1_40/Y vdd NAND3X1
XNAND3X1_73 NAND2X1_42/Y OR2X2_2/Y NAND2X1_41/Y gnd NAND3X1_74/A vdd NAND3X1
XNAND3X1_51 NAND3X1_44/Y NAND3X1_51/B NAND3X1_47/Y gnd OR2X2_2/A vdd NAND3X1
XNOR2X1_40 NOR2X1_40/A NOR2X1_40/B gnd NOR2X1_40/Y vdd NOR2X1
XNAND2X1_6 INVX1_2/A INVX2_1/A gnd INVX2_2/A vdd NAND2X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_21 NOR3X1_1/B gnd INVX1_21/Y vdd INVX1
XDFFPOSX1_6 DFFPOSX1_6/Q CLKBUF1_1/Y D[0] gnd vdd DFFPOSX1
XXNOR2X1_19 C[2] D[2] gnd XOR2X1_13/B vdd XNOR2X1
XINVX1_32 C[2] gnd INVX1_32/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd INVX2_5/A vdd NOR2X1
XAOI21X1_19 NAND3X1_28/Y NAND3X1_29/Y INVX2_5/Y gnd NOR3X1_2/A vdd AOI21X1
XOAI21X1_60 NOR2X1_4/A NOR2X1_1/B NOR2X1_3/B gnd AND2X2_10/B vdd OAI21X1
XFILL_8_1 gnd vdd FILL
XDFFPOSX1_19 NAND2X1_34/A CLKBUF1_6/Y DFFPOSX1_11/Q gnd vdd DFFPOSX1
XFILL_6_1_0 gnd vdd FILL
XNAND3X1_63 INVX1_18/Y NAND3X1_61/Y NAND3X1_62/Y gnd NAND3X1_63/Y vdd NAND3X1
XNOR2X1_41 NOR2X1_40/Y INVX1_46/Y gnd NOR2X1_41/Y vdd NOR2X1
XNAND3X1_41 OAI21X1_40/B OAI21X1_40/C AOI21X1_39/B gnd NAND3X1_46/A vdd NAND3X1
XNAND3X1_30 NOR3X1_1/Y NAND3X1_72/B OAI21X1_21/Y gnd XNOR2X1_3/B vdd NAND3X1
XNOR2X1_30 C[0] INVX1_30/Y gnd NOR2X1_30/Y vdd NOR2X1
XNAND3X1_74 NAND3X1_74/A AOI21X1_49/Y OAI21X1_46/Y gnd NAND2X1_43/A vdd NAND3X1
XNAND3X1_52 NAND3X1_49/Y NAND3X1_48/C OAI21X1_33/Y gnd AOI22X1_6/D vdd NAND3X1
XNAND2X1_7 BUFX4_7/Y AOI22X1_3/B gnd NOR2X1_5/B vdd NAND2X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_22 B[1] gnd INVX1_22/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_33 C[3] gnd INVX1_33/Y vdd INVX1
XDFFPOSX1_7 DFFPOSX1_7/Q CLKBUF1_1/Y D[1] gnd vdd DFFPOSX1
XOAI21X1_61 NOR2X1_8/Y NOR3X1_1/B NOR3X1_1/A gnd AND2X2_11/B vdd OAI21X1
XOAI21X1_50 C[0] INVX1_30/Y XNOR2X1_18/A gnd OAI21X1_51/C vdd OAI21X1
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_20 B[2] A[2] gnd NOR2X1_20/Y vdd NOR2X1
XNAND3X1_64 INVX1_19/A AOI21X1_46/A AOI21X1_46/B gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_42 AOI21X1_39/A NAND3X1_39/B NAND3X1_37/Y gnd NAND3X1_42/Y vdd NAND3X1
XNAND3X1_31 BUFX4_6/Y AOI22X1_5/B NOR2X1_13/A gnd NAND3X1_33/B vdd NAND3X1
XNAND3X1_75 INVX1_45/A INVX1_48/Y INVX1_46/A gnd AND2X2_8/B vdd NAND3X1
XNOR2X1_31 D[4] INVX1_34/Y gnd INVX1_35/A vdd NOR2X1
XNAND3X1_53 OR2X2_2/A AOI22X1_6/D NOR3X1_2/Y gnd NAND3X1_53/Y vdd NAND3X1
XNOR2X1_42 NOR2X1_42/A NOR2X1_42/B gnd NOR2X1_42/Y vdd NOR2X1
XNAND3X1_20 OAI22X1_2/Y NAND3X1_15/Y OAI21X1_18/Y gnd NAND3X1_20/Y vdd NAND3X1
XNAND2X1_8 INVX2_2/Y NOR2X1_6/Y gnd NAND3X1_1/C vdd NAND2X1
XINVX1_23 A[1] gnd INVX1_23/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_34 C[4] gnd INVX1_34/Y vdd INVX1
XDFFPOSX1_8 DFFPOSX1_8/Q CLKBUF1_5/Y D[2] gnd vdd DFFPOSX1
XOAI21X1_40 AOI21X1_42/Y OAI21X1_40/B OAI21X1_40/C gnd AOI21X1_43/C vdd OAI21X1
XOAI21X1_51 INVX1_31/Y D[1] OAI21X1_51/C gnd XOR2X1_13/A vdd OAI21X1
XAND2X2_10 INVX1_50/Y AND2X2_10/B gnd AND2X2_10/Y vdd AND2X2
XNAND3X1_65 INVX1_19/Y AOI21X1_45/A AOI21X1_45/B gnd NAND3X1_66/B vdd NAND3X1
XNOR2X1_21 NOR2X1_20/Y AND2X2_3/Y gnd XOR2X1_7/B vdd NOR2X1
XNAND3X1_32 BUFX4_2/Y INVX1_15/A NOR2X1_13/B gnd NAND3X1_32/Y vdd NAND3X1
XNAND3X1_54 NAND3X1_54/A BUFX4_5/Y OAI22X1_5/B gnd AOI21X1_37/A vdd NAND3X1
XNAND3X1_43 NAND3X1_46/A NAND3X1_45/B NAND3X1_42/Y gnd AOI21X1_33/B vdd NAND3X1
XNOR2X1_10 INVX1_11/Y INVX4_1/Y gnd XOR2X1_1/B vdd NOR2X1
XNOR2X1_43 NOR2X1_42/Y INVX1_47/Y gnd INVX1_48/A vdd NOR2X1
XNAND3X1_10 INVX1_10/Y NAND3X1_9/Y NAND3X1_8/Y gnd NAND3X1_10/Y vdd NAND3X1
XNAND3X1_21 OAI21X1_23/B NAND3X1_19/Y NAND3X1_20/Y gnd NAND3X1_21/Y vdd NAND3X1
XNOR2X1_32 INVX1_37/Y INVX2_8/Y gnd NOR2X1_32/Y vdd NOR2X1
XNAND2X1_9 INVX1_7/A INVX2_1/A gnd NAND3X1_8/C vdd NAND2X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 B[3] gnd INVX1_24/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XDFFPOSX1_9 DFFPOSX1_9/Q CLKBUF1_2/Y D[3] gnd vdd DFFPOSX1
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_41 OAI21X1_41/A OAI21X1_41/B INVX1_18/A gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_30 OAI21X1_30/A OAI21X1_30/B INVX1_12/Y gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_52 INVX1_32/Y D[2] NAND2X1_49/Y gnd XOR2X1_14/A vdd OAI21X1
XAND2X2_11 AND2X2_11/A AND2X2_11/B gnd AND2X2_11/Y vdd AND2X2
XFILL_6_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XNAND3X1_66 NAND3X1_64/Y NAND3X1_66/B NAND3X1_66/C gnd NAND3X1_66/Y vdd NAND3X1
XNAND3X1_33 INVX1_13/A NAND3X1_33/B NAND3X1_32/Y gnd NAND3X1_37/B vdd NAND3X1
XNAND3X1_55 BUFX4_1/Y AOI22X1_5/B NAND2X1_38/Y gnd AOI21X1_37/B vdd NAND3X1
XNOR2X1_22 INVX1_24/Y INVX1_25/Y gnd INVX1_26/A vdd NOR2X1
XNOR2X1_11 OAI22X1_4/A XOR2X1_3/A gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_33 AND2X2_7/A AND2X2_7/B gnd NOR2X1_33/Y vdd NOR2X1
XNAND3X1_22 NAND3X1_17/Y NAND3X1_21/Y AOI21X1_18/C gnd OAI21X1_32/C vdd NAND3X1
XNOR2X1_44 INVX1_47/Y INVX1_49/A gnd XOR2X1_22/A vdd NOR2X1
XNAND3X1_44 XOR2X1_1/Y AOI21X1_33/B NAND3X1_40/Y gnd NAND3X1_44/Y vdd NAND3X1
XNAND3X1_11 BUFX4_6/Y INVX1_15/A NOR2X1_12/A gnd NAND3X1_11/Y vdd NAND3X1
XINVX1_25 A[3] gnd INVX1_25/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_36 C[5] gnd OR2X2_3/A vdd INVX1
XINVX1_14 BUFX4_7/Y gnd INVX1_14/Y vdd INVX1
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_31 NOR2X1_11/Y AOI22X1_3/Y INVX1_12/A gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_42 AOI21X1_31/Y XNOR2X1_2/Y NAND3X1_40/Y gnd AOI21X1_47/C vdd OAI21X1
XOAI21X1_20 AOI21X1_17/Y OAI21X1_32/A INVX2_5/Y gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_53 INVX1_33/Y D[3] NAND2X1_50/Y gnd XNOR2X1_21/A vdd OAI21X1
XFILL_1_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XNAND3X1_67 AOI21X1_47/C OAI21X1_43/Y NAND3X1_66/Y gnd NAND2X1_41/B vdd NAND3X1
XNAND3X1_34 OAI22X1_3/Y NAND3X1_37/B NAND3X1_37/C gnd OAI21X1_40/C vdd NAND3X1
XNAND3X1_56 INVX1_17/Y AOI21X1_37/A AOI21X1_37/B gnd AOI21X1_36/A vdd NAND3X1
XNAND3X1_45 NAND3X1_36/Y NAND3X1_45/B AOI21X1_31/B gnd NAND3X1_47/B vdd NAND3X1
XNOR2X1_12 NOR2X1_12/A OAI22X1_5/A gnd NOR2X1_12/Y vdd NOR2X1
XNAND3X1_23 OAI21X1_23/B OAI21X1_23/C NAND3X1_16/Y gnd NAND3X1_23/Y vdd NAND3X1
XNAND3X1_12 BUFX4_2/Y AOI22X1_4/D OAI22X1_5/A gnd NAND3X1_12/Y vdd NAND3X1
XNOR2X1_23 B[3] A[3] gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_45 AND2X2_6/A AND2X2_6/B gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_34 NOR2X1_33/Y AND2X2_7/Y gnd XOR2X1_20/B vdd NOR2X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XOAI21X1_43 AOI21X1_45/Y AOI21X1_46/Y XOR2X1_4/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_21 NOR3X1_2/A NOR3X1_2/C OR2X2_1/Y gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_32 OAI21X1_32/A INVX2_5/Y OAI21X1_32/C gnd NAND3X1_51/B vdd OAI21X1
XOAI21X1_10 NOR2X1_7/Y AOI22X1_2/Y INVX2_3/A gnd AOI21X1_9/A vdd OAI21X1
XOAI21X1_54 INVX1_37/Y INVX1_35/Y OR2X2_3/Y gnd AOI21X1_53/C vdd OAI21X1
XNAND3X1_57 AOI21X1_36/A AOI21X1_36/B INVX1_16/Y gnd NAND3X1_57/Y vdd NAND3X1
XNOR2X1_35 INVX1_42/Y INVX1_43/Y gnd NOR2X1_37/B vdd NOR2X1
XNOR2X1_24 NOR2X1_23/Y INVX1_26/A gnd NOR2X1_24/Y vdd NOR2X1
XNAND3X1_68 AOI21X1_33/Y NAND3X1_63/Y OAI21X1_41/Y gnd NAND2X1_41/A vdd NAND3X1
XNAND3X1_35 AOI21X1_38/C AOI21X1_38/A AOI21X1_38/B gnd AOI21X1_39/B vdd NAND3X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XNAND3X1_46 NAND3X1_46/A NAND3X1_42/Y AOI21X1_31/C gnd NAND3X1_47/C vdd NAND3X1
XNOR2X1_46 NOR2X1_45/Y AND2X2_6/Y gnd NOR2X1_46/Y vdd NOR2X1
XNAND3X1_24 AOI21X1_29/A NAND3X1_19/Y NAND3X1_20/Y gnd NAND3X1_24/Y vdd NAND3X1
XNAND3X1_13 INVX2_4/A NAND3X1_11/Y NAND3X1_12/Y gnd NAND3X1_14/B vdd NAND3X1
XINVX1_16 NOR3X1_4/A gnd INVX1_16/Y vdd INVX1
XINVX1_38 D[6] gnd INVX1_38/Y vdd INVX1
XINVX1_27 B[5] gnd INVX1_27/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XOAI21X1_55 XOR2X1_16/A XOR2X1_16/B NAND2X1_53/Y gnd XNOR2X1_23/A vdd OAI21X1
XOAI21X1_44 AND2X2_1/Y NOR2X1_18/Y NAND2X1_41/Y gnd NAND3X1_69/B vdd OAI21X1
XOAI21X1_22 NOR2X1_9/B AOI21X1_24/C NAND2X1_23/B gnd XOR2X1_1/A vdd OAI21X1
XOAI21X1_33 AOI21X1_33/C AOI21X1_31/Y XOR2X1_1/Y gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_11 AOI21X1_5/Y AOI21X1_6/Y INVX2_3/A gnd NAND3X1_6/C vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XNAND3X1_58 NAND3X1_58/A NAND3X1_57/Y XNOR2X1_7/Y gnd AOI21X1_45/A vdd NAND3X1
XNOR2X1_36 INVX1_42/A INVX1_43/A gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_36 AOI21X1_39/A OAI21X1_40/C AOI21X1_39/B gnd NAND3X1_36/Y vdd NAND3X1
XNOR2X1_47 NOR2X1_47/A INVX1_20/Y gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_14 NOR3X1_2/A NOR3X1_2/C gnd NOR2X1_14/Y vdd NOR2X1
XNAND3X1_69 OAI21X1_34/Y NAND3X1_69/B NAND2X1_40/Y gnd NAND2X1_43/B vdd NAND3X1
XNAND3X1_25 NAND3X1_23/Y NAND3X1_24/Y NAND3X1_28/C gnd NAND3X1_25/Y vdd NAND3X1
XNOR2X1_25 INVX1_27/Y INVX1_28/Y gnd NOR2X1_25/Y vdd NOR2X1
XNAND3X1_14 OAI22X1_2/Y NAND3X1_14/B OAI21X1_17/Y gnd OAI21X1_23/C vdd NAND3X1
XNAND3X1_47 XNOR2X1_2/Y NAND3X1_47/B NAND3X1_47/C gnd NAND3X1_47/Y vdd NAND3X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_28 A[5] gnd INVX1_28/Y vdd INVX1
XOAI21X1_34 AOI22X1_6/Y XNOR2X1_3/B NAND3X1_53/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 NOR3X1_2/A NOR3X1_2/C NOR2X1_8/Y gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_12 NOR2X1_7/Y AOI22X1_2/Y INVX2_3/Y gnd NAND3X1_6/A vdd OAI21X1
XOAI21X1_23 AOI21X1_22/Y OAI21X1_23/B OAI21X1_23/C gnd AOI21X1_31/C vdd OAI21X1
XOAI21X1_56 INVX1_39/Y INVX1_40/Y NAND2X1_54/Y gnd XOR2X1_20/A vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XFILL_4_2 gnd vdd FILL
XNAND3X1_59 XOR2X1_3/Y AOI21X1_36/A AOI21X1_36/B gnd NAND3X1_59/Y vdd NAND3X1
XNOR2X1_37 NOR2X1_36/Y NOR2X1_37/B gnd INVX1_44/A vdd NOR2X1
XNAND3X1_37 AOI21X1_38/C NAND3X1_37/B NAND3X1_37/C gnd NAND3X1_37/Y vdd NAND3X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_15 NOR2X1_15/A AOI22X1_6/Y gnd XNOR2X1_3/A vdd NOR2X1
XNAND3X1_26 INVX2_5/A NAND3X1_25/Y OAI21X1_32/C gnd NAND3X1_27/B vdd NAND3X1
XNOR2X1_26 B[5] A[5] gnd INVX1_29/A vdd NOR2X1
XNAND3X1_48 NAND3X1_44/Y NAND3X1_47/Y NAND3X1_48/C gnd NAND3X1_48/Y vdd NAND3X1
XNAND3X1_15 INVX2_4/Y NAND3X1_11/Y NAND3X1_12/Y gnd NAND3X1_15/Y vdd NAND3X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XOAI21X1_35 NOR3X1_3/A NOR3X1_3/C INVX1_17/A gnd AOI21X1_36/B vdd OAI21X1
XOAI21X1_57 XNOR2X1_24/A INVX1_41/Y NAND2X1_55/Y gnd XNOR2X1_25/A vdd OAI21X1
XOAI21X1_24 OAI21X1_30/A OAI21X1_30/B INVX1_12/A gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_46 AND2X2_1/Y NOR2X1_18/Y NOR2X1_17/Y gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_13 AOI21X1_8/Y AOI21X1_9/Y INVX1_8/A gnd OAI21X1_13/Y vdd OAI21X1
XNAND3X1_38 OAI22X1_3/Y AOI21X1_38/A AOI21X1_38/B gnd NAND3X1_39/B vdd NAND3X1
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNAND3X1_27 NOR2X1_8/Y NAND3X1_27/B OAI21X1_20/Y gnd NAND3X1_72/B vdd NAND3X1
XNOR2X1_16 INVX1_11/Y INVX2_1/Y gnd XOR2X1_2/B vdd NOR2X1
XNOR2X1_27 INVX1_29/A NOR2X1_25/Y gnd NOR2X1_27/Y vdd NOR2X1
XNAND3X1_16 NAND3X1_19/A NAND3X1_15/Y OAI21X1_18/Y gnd NAND3X1_16/Y vdd NAND3X1
XNAND3X1_49 XNOR2X1_2/Y AOI21X1_33/B NAND3X1_40/Y gnd NAND3X1_49/Y vdd NAND3X1
XFILL_10_0_0 gnd vdd FILL
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_36 NOR3X1_4/Y AOI21X1_36/Y XNOR2X1_6/Y gnd AOI21X1_45/B vdd OAI21X1
XOAI21X1_47 INVX1_22/Y INVX1_23/Y OAI21X1_47/C gnd XOR2X1_7/A vdd OAI21X1
XOAI21X1_58 INVX1_42/Y INVX1_43/Y OAI21X1_58/C gnd NOR2X1_40/B vdd OAI21X1
XOAI21X1_25 NOR2X1_11/Y AOI22X1_3/Y INVX1_12/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_14 OAI21X1_6/B INVX1_5/A NAND3X1_3/B gnd OAI21X1_14/Y vdd OAI21X1
XXNOR2X1_1 XNOR2X1_1/A INVX1_3/Y gnd NOR2X1_3/B vdd XNOR2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_2_1 gnd vdd FILL
XAND2X2_1 OR2X2_2/A INVX2_7/Y gnd AND2X2_1/Y vdd AND2X2
XNOR2X1_17 NOR2X1_17/A NOR2X1_17/B gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_28 B[0] A[0] gnd NOR2X1_29/A vdd NOR2X1
XNAND3X1_39 OAI21X1_40/B NAND3X1_39/B NAND3X1_37/Y gnd AOI21X1_31/B vdd NAND3X1
XNAND3X1_28 NAND3X1_17/Y NAND3X1_21/Y NAND3X1_28/C gnd NAND3X1_28/Y vdd NAND3X1
XNAND3X1_17 AOI21X1_29/A OAI21X1_23/C NAND3X1_16/Y gnd NAND3X1_17/Y vdd NAND3X1
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_39 NOR2X1_38/Y INVX1_45/Y gnd NOR2X1_40/A vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XNAND2X1_50 XOR2X1_14/B XOR2X1_14/A gnd NAND2X1_50/Y vdd NAND2X1
XOAI21X1_37 NOR3X1_4/C NOR3X1_4/B NOR3X1_4/A gnd NAND3X1_58/A vdd OAI21X1
XOAI21X1_48 AOI21X1_50/Y NOR2X1_23/Y INVX1_26/Y gnd XOR2X1_9/A vdd OAI21X1
XOAI21X1_26 OAI21X1_26/A OAI21X1_26/B INVX1_13/Y gnd NAND3X1_37/C vdd OAI21X1
XOAI21X1_59 INVX1_4/Y INVX4_1/Y NOR2X1_4/A gnd AND2X2_9/B vdd OAI21X1
XOAI21X1_15 AOI21X1_9/Y INVX1_8/A NAND3X1_7/B gnd AOI21X1_18/C vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XXNOR2X1_2 XOR2X1_1/A XOR2X1_1/B gnd XNOR2X1_2/Y vdd XNOR2X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XAND2X2_2 B[0] A[0] gnd AND2X2_2/Y vdd AND2X2
XFILL_2_2 gnd vdd FILL
XNOR2X1_29 NOR2X1_29/A AND2X2_2/Y gnd NOR2X1_29/Y vdd NOR2X1
XNOR2X1_18 INVX2_7/Y OR2X2_2/A gnd NOR2X1_18/Y vdd NOR2X1
XNAND3X1_29 NAND3X1_23/Y NAND3X1_24/Y AOI21X1_18/C gnd NAND3X1_29/Y vdd NAND3X1
XNAND3X1_18 INVX1_10/A NAND3X1_9/Y NAND3X1_8/Y gnd NAND3X1_18/Y vdd NAND3X1
XNAND2X1_51 D[4] INVX1_34/Y gnd AND2X2_4/B vdd NAND2X1
XNAND2X1_40 NOR2X1_17/Y NAND2X1_40/B gnd NAND2X1_40/Y vdd NAND2X1
XOAI21X1_38 NOR3X1_4/C NOR3X1_4/B NOR3X1_5/A gnd NAND3X1_60/C vdd OAI21X1
XOAI21X1_49 XOR2X1_11/A XOR2X1_11/B NAND2X1_48/Y gnd XNOR2X1_16/A vdd OAI21X1
XOAI21X1_16 AOI21X1_11/Y OAI21X1_16/B INVX1_10/A gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_27 INVX1_14/Y INVX1_15/Y NOR2X1_12/A gnd OAI21X1_27/Y vdd OAI21X1
XXNOR2X1_3 XNOR2X1_3/A XNOR2X1_3/B gnd XNOR2X1_3/Y vdd XNOR2X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 B[2] A[2] gnd AND2X2_3/Y vdd AND2X2
XNOR2X1_19 INVX1_14/Y INVX4_1/Y gnd NOR2X1_19/Y vdd NOR2X1
XNAND3X1_19 NAND3X1_19/A NAND3X1_14/B OAI21X1_17/Y gnd NAND3X1_19/Y vdd NAND3X1
XNAND2X1_30 INVX1_2/A AOI22X1_4/D gnd INVX1_13/A vdd NAND2X1
XNAND2X1_41 NAND2X1_41/A NAND2X1_41/B gnd NAND2X1_41/Y vdd NAND2X1
XNAND2X1_52 D[5] OR2X2_3/A gnd AND2X2_5/B vdd NAND2X1
XOAI22X1_1 OAI22X1_1/A NOR2X1_7/A INVX1_9/A INVX2_2/A gnd NAND3X1_5/A vdd OAI22X1
XOAI21X1_39 NOR3X1_5/Y AOI21X1_41/Y XNOR2X1_9/Y gnd AOI21X1_46/B vdd OAI21X1
XOAI21X1_28 OAI21X1_26/A OAI21X1_26/B INVX1_13/A gnd AOI21X1_38/B vdd OAI21X1
XOAI21X1_17 OAI21X1_17/A OAI21X1_17/B INVX2_4/Y gnd OAI21X1_17/Y vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XXNOR2X1_4 XOR2X1_2/Y XNOR2X1_4/B gnd INVX1_18/A vdd XNOR2X1
XOR2X2_2 OR2X2_2/A INVX2_7/Y gnd OR2X2_2/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XAND2X2_4 INVX1_35/Y AND2X2_4/B gnd INVX2_8/A vdd AND2X2
XNAND2X1_31 BUFX4_8/Y AOI22X1_5/B gnd NOR2X1_13/B vdd NAND2X1
XNAND2X1_53 C[6] INVX1_38/Y gnd NAND2X1_53/Y vdd NAND2X1
XNAND2X1_42 INVX2_7/Y OR2X2_2/A gnd NAND2X1_42/Y vdd NAND2X1
XNAND2X1_20 INVX1_2/A AOI22X1_3/B gnd INVX2_4/A vdd NAND2X1
XOAI22X1_2 NOR2X1_5/B NOR2X1_12/A AOI22X1_2/Y INVX2_3/A gnd OAI22X1_2/Y vdd OAI22X1
XOAI21X1_29 NOR2X1_13/Y OAI22X1_5/C INVX1_13/Y gnd AOI21X1_38/A vdd OAI21X1
XOAI21X1_18 OAI21X1_17/A OAI21X1_17/B INVX2_4/A gnd OAI21X1_18/Y vdd OAI21X1
XFILL_12_2 gnd vdd FILL
XXNOR2X1_5 XOR2X1_3/A XOR2X1_3/B gnd NOR3X1_5/A vdd XNOR2X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOR2X2_3 OR2X2_3/A D[5] gnd OR2X2_3/Y vdd OR2X2
.ends

